module Multiplier 
import types::*;
(
    input clk,
    input rst,
    input logic mul_en,
    input logic [31:0] multiplier,
    input logic [31:0] multiplicand,
    input m_funct3_t mul_funct3,
    output logic [31:0] mul_out,
    output logic resp
);

logic [31:0] A, B;
logic [63:0] pre_result, pre_result_in;
logic [63:0] result;
// sign = 0 if both A and B are + or -; 
// sign = 1 if either is -; 
logic sign, sign_in; 

enum int unsigned {IDLE, PREPARE, REDUCTION} state, next_state;

always_ff @(posedge clk) begin
    if(rst) begin
        state <= IDLE;
        pre_result <= '0;
        sign <= 1'b0;
    end
    else begin
        state <= next_state;
        pre_result <= pre_result_in;
        sign <= sign_in;
    end
end

always_comb begin
    next_state = state;
    unique case (state)
        IDLE: begin
            if(mul_en)
                next_state = PREPARE;
            else 
                next_state = IDLE;
        end
        PREPARE: next_state = REDUCTION;
        REDUCTION: next_state = IDLE;
        default:;
    endcase
end

always_comb begin
    mul_out = 32'd0;
    resp = 1'b0;
    mul_out = '0;
    result = '0;
    sign_in = 1'b0;
    A = '0;
    B = '0;
    unique case (state)
        IDLE: begin 
            sign_in = 1'b0;
        end
        PREPARE:begin
            case (mul_funct3)
                mul, mulh: begin
                    if (multiplier[31] && !multiplicand[31]) begin      // A is -
                        sign_in = 1'b1;
                        A = ~multiplier + 1;
                        B = multiplicand;
                    end
                    else if(!multiplier[31] && multiplicand[31]) begin  // B is -
                        sign_in = 1'b1;
                        A = multiplier;
                        B = ~multiplicand + 1;
                    end
                    else if (multiplier[31] && multiplicand[31])begin   // A and B both -
                        sign_in = 1'b0;
                        A = ~multiplier + 1;
                        B = ~multiplicand + 1;
                    end
                    else begin                                          // A and B both +
                        sign_in = 1'b0;
                        A = multiplier;
                        B = multiplicand;
                    end
                end
                mulhsu: begin
                    if (multiplier[31]) begin      // A is -
                        sign_in = 1'b1;
                        A = ~multiplier + 1;
                        B = multiplicand;
                    end
                    else begin
                        sign_in = 1'b0;
                        A = multiplier;
                        B = multiplicand;
                    end
                end
                mulhu: begin
                    sign_in = 1'b0;
                    A = multiplier;
                    B = multiplicand;
                end
                default: begin
                    sign_in = 1'b0;
                    A = multiplier;
                    B = multiplicand;
                end
            endcase
        end
        REDUCTION: begin
            case (sign) 
                1'b0: result = pre_result;
                1'b1: result = ~pre_result + 1;
                default: result = '0;
            endcase
            case (mul_funct3) 
                mul: begin
                    mul_out = result[31:0];
                end
                default: begin
                    mul_out = result[63:32];
                end
            endcase
            resp = 1'b1;
        end
        default: begin
            sign_in = 1'b0;
            resp = 1'b0;
            mul_out = '0;
            result = '0;
            A = '0;
            B = '0;
        end
    endcase
end

logic ps_00, ps_11, ps_10, ps_22, ps_21, ps_20, ps_33, ps_32, ps_31, ps_30, ps_44, ps_43, ps_42, ps_41, ps_40, ps_55, ps_54, ps_53, ps_52, ps_51, ps_50, ps_66, ps_65, ps_64, ps_63, ps_62, ps_61, ps_60, ps_77, ps_76, ps_75, ps_74, ps_73, ps_72, ps_71, ps_70, ps_88, ps_87, ps_86, ps_85, ps_84, ps_83, ps_82, ps_81, ps_80, ps_99, ps_98, ps_97, ps_96, ps_95, ps_94, ps_93, ps_92, ps_91, ps_90, ps_1010, ps_109, ps_108, ps_107, ps_106, ps_105, ps_104, ps_103, ps_102, ps_101, ps_100, ps_1111, ps_1110, ps_119, ps_118, ps_117, ps_116, ps_115, ps_114, ps_113, ps_112, ps_111, ps_110, ps_1212, ps_1211, ps_1210, ps_129, ps_128, ps_127, ps_126, ps_125, ps_124, ps_123, ps_122, ps_121, ps_120, ps_1313, ps_1312, ps_1311, ps_1310, ps_139, ps_138, ps_137, ps_136, ps_135, ps_134, ps_133, ps_132, ps_131, ps_130, ps_1414, ps_1413, ps_1412, ps_1411, ps_1410, ps_149, ps_148, ps_147, ps_146, ps_145, ps_144, ps_143, ps_142, ps_141, ps_140, ps_1515, ps_1514, ps_1513, ps_1512, ps_1511, ps_1510, ps_159, ps_158, ps_157, ps_156, ps_155, ps_154, ps_153, ps_152, ps_151, ps_150, ps_1616, ps_1615, ps_1614, ps_1613, ps_1612, ps_1611, ps_1610, ps_169, ps_168, ps_167, ps_166, ps_165, ps_164, ps_163, ps_162, ps_161, ps_160, ps_1717, ps_1716, ps_1715, ps_1714, ps_1713, ps_1712, ps_1711, ps_1710, ps_179, ps_178, ps_177, ps_176, ps_175, ps_174, ps_173, ps_172, ps_171, ps_170, ps_1818, ps_1817, ps_1816, ps_1815, ps_1814, ps_1813, ps_1812, ps_1811, ps_1810, ps_189, ps_188, ps_187, ps_186, ps_185, ps_184, ps_183, ps_182, ps_181, ps_180, ps_1919, ps_1918, ps_1917, ps_1916, ps_1915, ps_1914, ps_1913, ps_1912, ps_1911, ps_1910, ps_199, ps_198, ps_197, ps_196, ps_195, ps_194, ps_193, ps_192, ps_191, ps_190, ps_2020, ps_2019, ps_2018, ps_2017, ps_2016, ps_2015, ps_2014, ps_2013, ps_2012, ps_2011, ps_2010, ps_209, ps_208, ps_207, ps_206, ps_205, ps_204, ps_203, ps_202, ps_201, ps_200, ps_2121, ps_2120, ps_2119, ps_2118, ps_2117, ps_2116, ps_2115, ps_2114, ps_2113, ps_2112, ps_2111, ps_2110, ps_219, ps_218, ps_217, ps_216, ps_215, ps_214, ps_213, ps_212, ps_211, ps_210, ps_2222, ps_2221, ps_2220, ps_2219, ps_2218, ps_2217, ps_2216, ps_2215, ps_2214, ps_2213, ps_2212, ps_2211, ps_2210, ps_229, ps_228, ps_227, ps_226, ps_225, ps_224, ps_223, ps_222, ps_221, ps_220, ps_2323, ps_2322, ps_2321, ps_2320, ps_2319, ps_2318, ps_2317, ps_2316, ps_2315, ps_2314, ps_2313, ps_2312, ps_2311, ps_2310, ps_239, ps_238, ps_237, ps_236, ps_235, ps_234, ps_233, ps_232, ps_231, ps_230, ps_2424, ps_2423, ps_2422, ps_2421, ps_2420, ps_2419, ps_2418, ps_2417, ps_2416, ps_2415, ps_2414, ps_2413, ps_2412, ps_2411, ps_2410, ps_249, ps_248, ps_247, ps_246, ps_245, ps_244, ps_243, ps_242, ps_241, ps_240, ps_2525, ps_2524, ps_2523, ps_2522, ps_2521, ps_2520, ps_2519, ps_2518, ps_2517, ps_2516, ps_2515, ps_2514, ps_2513, ps_2512, ps_2511, ps_2510, ps_259, ps_258, ps_257, ps_256, ps_255, ps_254, ps_253, ps_252, ps_251, ps_250, ps_2626, ps_2625, ps_2624, ps_2623, ps_2622, ps_2621, ps_2620, ps_2619, ps_2618, ps_2617, ps_2616, ps_2615, ps_2614, ps_2613, ps_2612, ps_2611, ps_2610, ps_269, ps_268, ps_267, ps_266, ps_265, ps_264, ps_263, ps_262, ps_261, ps_260, ps_2727, ps_2726, ps_2725, ps_2724, ps_2723, ps_2722, ps_2721, ps_2720, ps_2719, ps_2718, ps_2717, ps_2716, ps_2715, ps_2714, ps_2713, ps_2712, ps_2711, ps_2710, ps_279, ps_278, ps_277, ps_276, ps_275, ps_274, ps_273, ps_272, ps_271, ps_270, ps_2828, ps_2827, ps_2826, ps_2825, ps_2824, ps_2823, ps_2822, ps_2821, ps_2820, ps_2819, ps_2818, ps_2817, ps_2816, ps_2815, ps_2814, ps_2813, ps_2812, ps_2811, ps_2810, ps_289, ps_288, ps_287, ps_286, ps_285, ps_284, ps_283, ps_282, ps_281, ps_280, ps_2929, ps_2928, ps_2927, ps_2926, ps_2925, ps_2924, ps_2923, ps_2922, ps_2921, ps_2920, ps_2919, ps_2918, ps_2917, ps_2916, ps_2915, ps_2914, ps_2913, ps_2912, ps_2911, ps_2910, ps_299, ps_298, ps_297, ps_296, ps_295, ps_294, ps_293, ps_292, ps_291, ps_290, ps_3030, ps_3029, ps_3028, ps_3027, ps_3026, ps_3025, ps_3024, ps_3023, ps_3022, ps_3021, ps_3020, ps_3019, ps_3018, ps_3017, ps_3016, ps_3015, ps_3014, ps_3013, ps_3012, ps_3011, ps_3010, ps_309, ps_308, ps_307, ps_306, ps_305, ps_304, ps_303, ps_302, ps_301, ps_300, ps_3131, ps_3130, ps_3129, ps_3128, ps_3127, ps_3126, ps_3125, ps_3124, ps_3123, ps_3122, ps_3121, ps_3120, ps_3119, ps_3118, ps_3117, ps_3116, ps_3115, ps_3114, ps_3113, ps_3112, ps_3111, ps_3110, ps_319, ps_318, ps_317, ps_316, ps_315, ps_314, ps_313, ps_312, ps_311, ps_310, ps_3231, ps_3230, ps_3229, ps_3228, ps_3227, ps_3226, ps_3225, ps_3224, ps_3223, ps_3222, ps_3221, ps_3220, ps_3219, ps_3218, ps_3217, ps_3216, ps_3215, ps_3214, ps_3213, ps_3212, ps_3211, ps_3210, ps_329, ps_328, ps_327, ps_326, ps_325, ps_324, ps_323, ps_322, ps_321, ps_3331, ps_3330, ps_3329, ps_3328, ps_3327, ps_3326, ps_3325, ps_3324, ps_3323, ps_3322, ps_3321, ps_3320, ps_3319, ps_3318, ps_3317, ps_3316, ps_3315, ps_3314, ps_3313, ps_3312, ps_3311, ps_3310, ps_339, ps_338, ps_337, ps_336, ps_335, ps_334, ps_333, ps_332, ps_3431, ps_3430, ps_3429, ps_3428, ps_3427, ps_3426, ps_3425, ps_3424, ps_3423, ps_3422, ps_3421, ps_3420, ps_3419, ps_3418, ps_3417, ps_3416, ps_3415, ps_3414, ps_3413, ps_3412, ps_3411, ps_3410, ps_349, ps_348, ps_347, ps_346, ps_345, ps_344, ps_343, ps_3531, ps_3530, ps_3529, ps_3528, ps_3527, ps_3526, ps_3525, ps_3524, ps_3523, ps_3522, ps_3521, ps_3520, ps_3519, ps_3518, ps_3517, ps_3516, ps_3515, ps_3514, ps_3513, ps_3512, ps_3511, ps_3510, ps_359, ps_358, ps_357, ps_356, ps_355, ps_354, ps_3631, ps_3630, ps_3629, ps_3628, ps_3627, ps_3626, ps_3625, ps_3624, ps_3623, ps_3622, ps_3621, ps_3620, ps_3619, ps_3618, ps_3617, ps_3616, ps_3615, ps_3614, ps_3613, ps_3612, ps_3611, ps_3610, ps_369, ps_368, ps_367, ps_366, ps_365, ps_3731, ps_3730, ps_3729, ps_3728, ps_3727, ps_3726, ps_3725, ps_3724, ps_3723, ps_3722, ps_3721, ps_3720, ps_3719, ps_3718, ps_3717, ps_3716, ps_3715, ps_3714, ps_3713, ps_3712, ps_3711, ps_3710, ps_379, ps_378, ps_377, ps_376, ps_3831, ps_3830, ps_3829, ps_3828, ps_3827, ps_3826, ps_3825, ps_3824, ps_3823, ps_3822, ps_3821, ps_3820, ps_3819, ps_3818, ps_3817, ps_3816, ps_3815, ps_3814, ps_3813, ps_3812, ps_3811, ps_3810, ps_389, ps_388, ps_387, ps_3931, ps_3930, ps_3929, ps_3928, ps_3927, ps_3926, ps_3925, ps_3924, ps_3923, ps_3922, ps_3921, ps_3920, ps_3919, ps_3918, ps_3917, ps_3916, ps_3915, ps_3914, ps_3913, ps_3912, ps_3911, ps_3910, ps_399, ps_398, ps_4031, ps_4030, ps_4029, ps_4028, ps_4027, ps_4026, ps_4025, ps_4024, ps_4023, ps_4022, ps_4021, ps_4020, ps_4019, ps_4018, ps_4017, ps_4016, ps_4015, ps_4014, ps_4013, ps_4012, ps_4011, ps_4010, ps_409, ps_4131, ps_4130, ps_4129, ps_4128, ps_4127, ps_4126, ps_4125, ps_4124, ps_4123, ps_4122, ps_4121, ps_4120, ps_4119, ps_4118, ps_4117, ps_4116, ps_4115, ps_4114, ps_4113, ps_4112, ps_4111, ps_4110, ps_4231, ps_4230, ps_4229, ps_4228, ps_4227, ps_4226, ps_4225, ps_4224, ps_4223, ps_4222, ps_4221, ps_4220, ps_4219, ps_4218, ps_4217, ps_4216, ps_4215, ps_4214, ps_4213, ps_4212, ps_4211, ps_4331, ps_4330, ps_4329, ps_4328, ps_4327, ps_4326, ps_4325, ps_4324, ps_4323, ps_4322, ps_4321, ps_4320, ps_4319, ps_4318, ps_4317, ps_4316, ps_4315, ps_4314, ps_4313, ps_4312, ps_4431, ps_4430, ps_4429, ps_4428, ps_4427, ps_4426, ps_4425, ps_4424, ps_4423, ps_4422, ps_4421, ps_4420, ps_4419, ps_4418, ps_4417, ps_4416, ps_4415, ps_4414, ps_4413, ps_4531, ps_4530, ps_4529, ps_4528, ps_4527, ps_4526, ps_4525, ps_4524, ps_4523, ps_4522, ps_4521, ps_4520, ps_4519, ps_4518, ps_4517, ps_4516, ps_4515, ps_4514, ps_4631, ps_4630, ps_4629, ps_4628, ps_4627, ps_4626, ps_4625, ps_4624, ps_4623, ps_4622, ps_4621, ps_4620, ps_4619, ps_4618, ps_4617, ps_4616, ps_4615, ps_4731, ps_4730, ps_4729, ps_4728, ps_4727, ps_4726, ps_4725, ps_4724, ps_4723, ps_4722, ps_4721, ps_4720, ps_4719, ps_4718, ps_4717, ps_4716, ps_4831, ps_4830, ps_4829, ps_4828, ps_4827, ps_4826, ps_4825, ps_4824, ps_4823, ps_4822, ps_4821, ps_4820, ps_4819, ps_4818, ps_4817, ps_4931, ps_4930, ps_4929, ps_4928, ps_4927, ps_4926, ps_4925, ps_4924, ps_4923, ps_4922, ps_4921, ps_4920, ps_4919, ps_4918, ps_5031, ps_5030, ps_5029, ps_5028, ps_5027, ps_5026, ps_5025, ps_5024, ps_5023, ps_5022, ps_5021, ps_5020, ps_5019, ps_5131, ps_5130, ps_5129, ps_5128, ps_5127, ps_5126, ps_5125, ps_5124, ps_5123, ps_5122, ps_5121, ps_5120, ps_5231, ps_5230, ps_5229, ps_5228, ps_5227, ps_5226, ps_5225, ps_5224, ps_5223, ps_5222, ps_5221, ps_5331, ps_5330, ps_5329, ps_5328, ps_5327, ps_5326, ps_5325, ps_5324, ps_5323, ps_5322, ps_5431, ps_5430, ps_5429, ps_5428, ps_5427, ps_5426, ps_5425, ps_5424, ps_5423, ps_5531, ps_5530, ps_5529, ps_5528, ps_5527, ps_5526, ps_5525, ps_5524, ps_5631, ps_5630, ps_5629, ps_5628, ps_5627, ps_5626, ps_5625, ps_5731, ps_5730, ps_5729, ps_5728, ps_5727, ps_5726, ps_5831, ps_5830, ps_5829, ps_5828, ps_5827, ps_5931, ps_5930, ps_5929, ps_5928, ps_6031, ps_6030, ps_6029, ps_6131, ps_6130, ps_6231;
assign ps_00 = A[0] & B[0]; 
assign ps_11 = A[1] & B[0]; 
assign ps_10 = A[0] & B[1]; 
assign ps_22 = A[2] & B[0]; 
assign ps_21 = A[1] & B[1]; 
assign ps_20 = A[0] & B[2]; 
assign ps_33 = A[3] & B[0]; 
assign ps_32 = A[2] & B[1]; 
assign ps_31 = A[1] & B[2]; 
assign ps_30 = A[0] & B[3]; 
assign ps_44 = A[4] & B[0]; 
assign ps_43 = A[3] & B[1]; 
assign ps_42 = A[2] & B[2]; 
assign ps_41 = A[1] & B[3]; 
assign ps_40 = A[0] & B[4]; 
assign ps_55 = A[5] & B[0]; 
assign ps_54 = A[4] & B[1]; 
assign ps_53 = A[3] & B[2]; 
assign ps_52 = A[2] & B[3]; 
assign ps_51 = A[1] & B[4]; 
assign ps_50 = A[0] & B[5]; 
assign ps_66 = A[6] & B[0]; 
assign ps_65 = A[5] & B[1]; 
assign ps_64 = A[4] & B[2]; 
assign ps_63 = A[3] & B[3]; 
assign ps_62 = A[2] & B[4]; 
assign ps_61 = A[1] & B[5]; 
assign ps_60 = A[0] & B[6]; 
assign ps_77 = A[7] & B[0]; 
assign ps_76 = A[6] & B[1]; 
assign ps_75 = A[5] & B[2]; 
assign ps_74 = A[4] & B[3]; 
assign ps_73 = A[3] & B[4]; 
assign ps_72 = A[2] & B[5]; 
assign ps_71 = A[1] & B[6]; 
assign ps_70 = A[0] & B[7]; 
assign ps_88 = A[8] & B[0]; 
assign ps_87 = A[7] & B[1]; 
assign ps_86 = A[6] & B[2]; 
assign ps_85 = A[5] & B[3]; 
assign ps_84 = A[4] & B[4]; 
assign ps_83 = A[3] & B[5]; 
assign ps_82 = A[2] & B[6]; 
assign ps_81 = A[1] & B[7]; 
assign ps_80 = A[0] & B[8]; 
assign ps_99 = A[9] & B[0]; 
assign ps_98 = A[8] & B[1]; 
assign ps_97 = A[7] & B[2]; 
assign ps_96 = A[6] & B[3]; 
assign ps_95 = A[5] & B[4]; 
assign ps_94 = A[4] & B[5]; 
assign ps_93 = A[3] & B[6]; 
assign ps_92 = A[2] & B[7]; 
assign ps_91 = A[1] & B[8]; 
assign ps_90 = A[0] & B[9]; 
assign ps_1010 = A[10] & B[0]; 
assign ps_109 = A[9] & B[1]; 
assign ps_108 = A[8] & B[2]; 
assign ps_107 = A[7] & B[3]; 
assign ps_106 = A[6] & B[4]; 
assign ps_105 = A[5] & B[5]; 
assign ps_104 = A[4] & B[6]; 
assign ps_103 = A[3] & B[7]; 
assign ps_102 = A[2] & B[8]; 
assign ps_101 = A[1] & B[9]; 
assign ps_100 = A[0] & B[10]; 
assign ps_1111 = A[11] & B[0]; 
assign ps_1110 = A[10] & B[1]; 
assign ps_119 = A[9] & B[2]; 
assign ps_118 = A[8] & B[3]; 
assign ps_117 = A[7] & B[4]; 
assign ps_116 = A[6] & B[5]; 
assign ps_115 = A[5] & B[6]; 
assign ps_114 = A[4] & B[7]; 
assign ps_113 = A[3] & B[8]; 
assign ps_112 = A[2] & B[9]; 
assign ps_111 = A[1] & B[10]; 
assign ps_110 = A[0] & B[11]; 
assign ps_1212 = A[12] & B[0]; 
assign ps_1211 = A[11] & B[1]; 
assign ps_1210 = A[10] & B[2]; 
assign ps_129 = A[9] & B[3]; 
assign ps_128 = A[8] & B[4]; 
assign ps_127 = A[7] & B[5]; 
assign ps_126 = A[6] & B[6]; 
assign ps_125 = A[5] & B[7]; 
assign ps_124 = A[4] & B[8]; 
assign ps_123 = A[3] & B[9]; 
assign ps_122 = A[2] & B[10]; 
assign ps_121 = A[1] & B[11]; 
assign ps_120 = A[0] & B[12]; 
assign ps_1313 = A[13] & B[0]; 
assign ps_1312 = A[12] & B[1]; 
assign ps_1311 = A[11] & B[2]; 
assign ps_1310 = A[10] & B[3]; 
assign ps_139 = A[9] & B[4]; 
assign ps_138 = A[8] & B[5]; 
assign ps_137 = A[7] & B[6]; 
assign ps_136 = A[6] & B[7]; 
assign ps_135 = A[5] & B[8]; 
assign ps_134 = A[4] & B[9]; 
assign ps_133 = A[3] & B[10]; 
assign ps_132 = A[2] & B[11]; 
assign ps_131 = A[1] & B[12]; 
assign ps_130 = A[0] & B[13]; 
assign ps_1414 = A[14] & B[0]; 
assign ps_1413 = A[13] & B[1]; 
assign ps_1412 = A[12] & B[2]; 
assign ps_1411 = A[11] & B[3]; 
assign ps_1410 = A[10] & B[4]; 
assign ps_149 = A[9] & B[5]; 
assign ps_148 = A[8] & B[6]; 
assign ps_147 = A[7] & B[7]; 
assign ps_146 = A[6] & B[8]; 
assign ps_145 = A[5] & B[9]; 
assign ps_144 = A[4] & B[10]; 
assign ps_143 = A[3] & B[11]; 
assign ps_142 = A[2] & B[12]; 
assign ps_141 = A[1] & B[13]; 
assign ps_140 = A[0] & B[14]; 
assign ps_1515 = A[15] & B[0]; 
assign ps_1514 = A[14] & B[1]; 
assign ps_1513 = A[13] & B[2]; 
assign ps_1512 = A[12] & B[3]; 
assign ps_1511 = A[11] & B[4]; 
assign ps_1510 = A[10] & B[5]; 
assign ps_159 = A[9] & B[6]; 
assign ps_158 = A[8] & B[7]; 
assign ps_157 = A[7] & B[8]; 
assign ps_156 = A[6] & B[9]; 
assign ps_155 = A[5] & B[10]; 
assign ps_154 = A[4] & B[11]; 
assign ps_153 = A[3] & B[12]; 
assign ps_152 = A[2] & B[13]; 
assign ps_151 = A[1] & B[14]; 
assign ps_150 = A[0] & B[15]; 
assign ps_1616 = A[16] & B[0]; 
assign ps_1615 = A[15] & B[1]; 
assign ps_1614 = A[14] & B[2]; 
assign ps_1613 = A[13] & B[3]; 
assign ps_1612 = A[12] & B[4]; 
assign ps_1611 = A[11] & B[5]; 
assign ps_1610 = A[10] & B[6]; 
assign ps_169 = A[9] & B[7]; 
assign ps_168 = A[8] & B[8]; 
assign ps_167 = A[7] & B[9]; 
assign ps_166 = A[6] & B[10]; 
assign ps_165 = A[5] & B[11]; 
assign ps_164 = A[4] & B[12]; 
assign ps_163 = A[3] & B[13]; 
assign ps_162 = A[2] & B[14]; 
assign ps_161 = A[1] & B[15]; 
assign ps_160 = A[0] & B[16]; 
assign ps_1717 = A[17] & B[0]; 
assign ps_1716 = A[16] & B[1]; 
assign ps_1715 = A[15] & B[2]; 
assign ps_1714 = A[14] & B[3]; 
assign ps_1713 = A[13] & B[4]; 
assign ps_1712 = A[12] & B[5]; 
assign ps_1711 = A[11] & B[6]; 
assign ps_1710 = A[10] & B[7]; 
assign ps_179 = A[9] & B[8]; 
assign ps_178 = A[8] & B[9]; 
assign ps_177 = A[7] & B[10]; 
assign ps_176 = A[6] & B[11]; 
assign ps_175 = A[5] & B[12]; 
assign ps_174 = A[4] & B[13]; 
assign ps_173 = A[3] & B[14]; 
assign ps_172 = A[2] & B[15]; 
assign ps_171 = A[1] & B[16]; 
assign ps_170 = A[0] & B[17]; 
assign ps_1818 = A[18] & B[0]; 
assign ps_1817 = A[17] & B[1]; 
assign ps_1816 = A[16] & B[2]; 
assign ps_1815 = A[15] & B[3]; 
assign ps_1814 = A[14] & B[4]; 
assign ps_1813 = A[13] & B[5]; 
assign ps_1812 = A[12] & B[6]; 
assign ps_1811 = A[11] & B[7]; 
assign ps_1810 = A[10] & B[8]; 
assign ps_189 = A[9] & B[9]; 
assign ps_188 = A[8] & B[10]; 
assign ps_187 = A[7] & B[11]; 
assign ps_186 = A[6] & B[12]; 
assign ps_185 = A[5] & B[13]; 
assign ps_184 = A[4] & B[14]; 
assign ps_183 = A[3] & B[15]; 
assign ps_182 = A[2] & B[16]; 
assign ps_181 = A[1] & B[17]; 
assign ps_180 = A[0] & B[18]; 
assign ps_1919 = A[19] & B[0]; 
assign ps_1918 = A[18] & B[1]; 
assign ps_1917 = A[17] & B[2]; 
assign ps_1916 = A[16] & B[3]; 
assign ps_1915 = A[15] & B[4]; 
assign ps_1914 = A[14] & B[5]; 
assign ps_1913 = A[13] & B[6]; 
assign ps_1912 = A[12] & B[7]; 
assign ps_1911 = A[11] & B[8]; 
assign ps_1910 = A[10] & B[9]; 
assign ps_199 = A[9] & B[10]; 
assign ps_198 = A[8] & B[11]; 
assign ps_197 = A[7] & B[12]; 
assign ps_196 = A[6] & B[13]; 
assign ps_195 = A[5] & B[14]; 
assign ps_194 = A[4] & B[15]; 
assign ps_193 = A[3] & B[16]; 
assign ps_192 = A[2] & B[17]; 
assign ps_191 = A[1] & B[18]; 
assign ps_190 = A[0] & B[19]; 
assign ps_2020 = A[20] & B[0]; 
assign ps_2019 = A[19] & B[1]; 
assign ps_2018 = A[18] & B[2]; 
assign ps_2017 = A[17] & B[3]; 
assign ps_2016 = A[16] & B[4]; 
assign ps_2015 = A[15] & B[5]; 
assign ps_2014 = A[14] & B[6]; 
assign ps_2013 = A[13] & B[7]; 
assign ps_2012 = A[12] & B[8]; 
assign ps_2011 = A[11] & B[9]; 
assign ps_2010 = A[10] & B[10]; 
assign ps_209 = A[9] & B[11]; 
assign ps_208 = A[8] & B[12]; 
assign ps_207 = A[7] & B[13]; 
assign ps_206 = A[6] & B[14]; 
assign ps_205 = A[5] & B[15]; 
assign ps_204 = A[4] & B[16]; 
assign ps_203 = A[3] & B[17]; 
assign ps_202 = A[2] & B[18]; 
assign ps_201 = A[1] & B[19]; 
assign ps_200 = A[0] & B[20]; 
assign ps_2121 = A[21] & B[0]; 
assign ps_2120 = A[20] & B[1]; 
assign ps_2119 = A[19] & B[2]; 
assign ps_2118 = A[18] & B[3]; 
assign ps_2117 = A[17] & B[4]; 
assign ps_2116 = A[16] & B[5]; 
assign ps_2115 = A[15] & B[6]; 
assign ps_2114 = A[14] & B[7]; 
assign ps_2113 = A[13] & B[8]; 
assign ps_2112 = A[12] & B[9]; 
assign ps_2111 = A[11] & B[10]; 
assign ps_2110 = A[10] & B[11]; 
assign ps_219 = A[9] & B[12]; 
assign ps_218 = A[8] & B[13]; 
assign ps_217 = A[7] & B[14]; 
assign ps_216 = A[6] & B[15]; 
assign ps_215 = A[5] & B[16]; 
assign ps_214 = A[4] & B[17]; 
assign ps_213 = A[3] & B[18]; 
assign ps_212 = A[2] & B[19]; 
assign ps_211 = A[1] & B[20]; 
assign ps_210 = A[0] & B[21]; 
assign ps_2222 = A[22] & B[0]; 
assign ps_2221 = A[21] & B[1]; 
assign ps_2220 = A[20] & B[2]; 
assign ps_2219 = A[19] & B[3]; 
assign ps_2218 = A[18] & B[4]; 
assign ps_2217 = A[17] & B[5]; 
assign ps_2216 = A[16] & B[6]; 
assign ps_2215 = A[15] & B[7]; 
assign ps_2214 = A[14] & B[8]; 
assign ps_2213 = A[13] & B[9]; 
assign ps_2212 = A[12] & B[10]; 
assign ps_2211 = A[11] & B[11]; 
assign ps_2210 = A[10] & B[12]; 
assign ps_229 = A[9] & B[13]; 
assign ps_228 = A[8] & B[14]; 
assign ps_227 = A[7] & B[15]; 
assign ps_226 = A[6] & B[16]; 
assign ps_225 = A[5] & B[17]; 
assign ps_224 = A[4] & B[18]; 
assign ps_223 = A[3] & B[19]; 
assign ps_222 = A[2] & B[20]; 
assign ps_221 = A[1] & B[21]; 
assign ps_220 = A[0] & B[22]; 
assign ps_2323 = A[23] & B[0]; 
assign ps_2322 = A[22] & B[1]; 
assign ps_2321 = A[21] & B[2]; 
assign ps_2320 = A[20] & B[3]; 
assign ps_2319 = A[19] & B[4]; 
assign ps_2318 = A[18] & B[5]; 
assign ps_2317 = A[17] & B[6]; 
assign ps_2316 = A[16] & B[7]; 
assign ps_2315 = A[15] & B[8]; 
assign ps_2314 = A[14] & B[9]; 
assign ps_2313 = A[13] & B[10]; 
assign ps_2312 = A[12] & B[11]; 
assign ps_2311 = A[11] & B[12]; 
assign ps_2310 = A[10] & B[13]; 
assign ps_239 = A[9] & B[14]; 
assign ps_238 = A[8] & B[15]; 
assign ps_237 = A[7] & B[16]; 
assign ps_236 = A[6] & B[17]; 
assign ps_235 = A[5] & B[18]; 
assign ps_234 = A[4] & B[19]; 
assign ps_233 = A[3] & B[20]; 
assign ps_232 = A[2] & B[21]; 
assign ps_231 = A[1] & B[22]; 
assign ps_230 = A[0] & B[23]; 
assign ps_2424 = A[24] & B[0]; 
assign ps_2423 = A[23] & B[1]; 
assign ps_2422 = A[22] & B[2]; 
assign ps_2421 = A[21] & B[3]; 
assign ps_2420 = A[20] & B[4]; 
assign ps_2419 = A[19] & B[5]; 
assign ps_2418 = A[18] & B[6]; 
assign ps_2417 = A[17] & B[7]; 
assign ps_2416 = A[16] & B[8]; 
assign ps_2415 = A[15] & B[9]; 
assign ps_2414 = A[14] & B[10]; 
assign ps_2413 = A[13] & B[11]; 
assign ps_2412 = A[12] & B[12]; 
assign ps_2411 = A[11] & B[13]; 
assign ps_2410 = A[10] & B[14]; 
assign ps_249 = A[9] & B[15]; 
assign ps_248 = A[8] & B[16]; 
assign ps_247 = A[7] & B[17]; 
assign ps_246 = A[6] & B[18]; 
assign ps_245 = A[5] & B[19]; 
assign ps_244 = A[4] & B[20]; 
assign ps_243 = A[3] & B[21]; 
assign ps_242 = A[2] & B[22]; 
assign ps_241 = A[1] & B[23]; 
assign ps_240 = A[0] & B[24]; 
assign ps_2525 = A[25] & B[0]; 
assign ps_2524 = A[24] & B[1]; 
assign ps_2523 = A[23] & B[2]; 
assign ps_2522 = A[22] & B[3]; 
assign ps_2521 = A[21] & B[4]; 
assign ps_2520 = A[20] & B[5]; 
assign ps_2519 = A[19] & B[6]; 
assign ps_2518 = A[18] & B[7]; 
assign ps_2517 = A[17] & B[8]; 
assign ps_2516 = A[16] & B[9]; 
assign ps_2515 = A[15] & B[10]; 
assign ps_2514 = A[14] & B[11]; 
assign ps_2513 = A[13] & B[12]; 
assign ps_2512 = A[12] & B[13]; 
assign ps_2511 = A[11] & B[14]; 
assign ps_2510 = A[10] & B[15]; 
assign ps_259 = A[9] & B[16]; 
assign ps_258 = A[8] & B[17]; 
assign ps_257 = A[7] & B[18]; 
assign ps_256 = A[6] & B[19]; 
assign ps_255 = A[5] & B[20]; 
assign ps_254 = A[4] & B[21]; 
assign ps_253 = A[3] & B[22]; 
assign ps_252 = A[2] & B[23]; 
assign ps_251 = A[1] & B[24]; 
assign ps_250 = A[0] & B[25]; 
assign ps_2626 = A[26] & B[0]; 
assign ps_2625 = A[25] & B[1]; 
assign ps_2624 = A[24] & B[2]; 
assign ps_2623 = A[23] & B[3]; 
assign ps_2622 = A[22] & B[4]; 
assign ps_2621 = A[21] & B[5]; 
assign ps_2620 = A[20] & B[6]; 
assign ps_2619 = A[19] & B[7]; 
assign ps_2618 = A[18] & B[8]; 
assign ps_2617 = A[17] & B[9]; 
assign ps_2616 = A[16] & B[10]; 
assign ps_2615 = A[15] & B[11]; 
assign ps_2614 = A[14] & B[12]; 
assign ps_2613 = A[13] & B[13]; 
assign ps_2612 = A[12] & B[14]; 
assign ps_2611 = A[11] & B[15]; 
assign ps_2610 = A[10] & B[16]; 
assign ps_269 = A[9] & B[17]; 
assign ps_268 = A[8] & B[18]; 
assign ps_267 = A[7] & B[19]; 
assign ps_266 = A[6] & B[20]; 
assign ps_265 = A[5] & B[21]; 
assign ps_264 = A[4] & B[22]; 
assign ps_263 = A[3] & B[23]; 
assign ps_262 = A[2] & B[24]; 
assign ps_261 = A[1] & B[25]; 
assign ps_260 = A[0] & B[26]; 
assign ps_2727 = A[27] & B[0]; 
assign ps_2726 = A[26] & B[1]; 
assign ps_2725 = A[25] & B[2]; 
assign ps_2724 = A[24] & B[3]; 
assign ps_2723 = A[23] & B[4]; 
assign ps_2722 = A[22] & B[5]; 
assign ps_2721 = A[21] & B[6]; 
assign ps_2720 = A[20] & B[7]; 
assign ps_2719 = A[19] & B[8]; 
assign ps_2718 = A[18] & B[9]; 
assign ps_2717 = A[17] & B[10]; 
assign ps_2716 = A[16] & B[11]; 
assign ps_2715 = A[15] & B[12]; 
assign ps_2714 = A[14] & B[13]; 
assign ps_2713 = A[13] & B[14]; 
assign ps_2712 = A[12] & B[15]; 
assign ps_2711 = A[11] & B[16]; 
assign ps_2710 = A[10] & B[17]; 
assign ps_279 = A[9] & B[18]; 
assign ps_278 = A[8] & B[19]; 
assign ps_277 = A[7] & B[20]; 
assign ps_276 = A[6] & B[21]; 
assign ps_275 = A[5] & B[22]; 
assign ps_274 = A[4] & B[23]; 
assign ps_273 = A[3] & B[24]; 
assign ps_272 = A[2] & B[25]; 
assign ps_271 = A[1] & B[26]; 
assign ps_270 = A[0] & B[27]; 
assign ps_2828 = A[28] & B[0]; 
assign ps_2827 = A[27] & B[1]; 
assign ps_2826 = A[26] & B[2]; 
assign ps_2825 = A[25] & B[3]; 
assign ps_2824 = A[24] & B[4]; 
assign ps_2823 = A[23] & B[5]; 
assign ps_2822 = A[22] & B[6]; 
assign ps_2821 = A[21] & B[7]; 
assign ps_2820 = A[20] & B[8]; 
assign ps_2819 = A[19] & B[9]; 
assign ps_2818 = A[18] & B[10]; 
assign ps_2817 = A[17] & B[11]; 
assign ps_2816 = A[16] & B[12]; 
assign ps_2815 = A[15] & B[13]; 
assign ps_2814 = A[14] & B[14]; 
assign ps_2813 = A[13] & B[15]; 
assign ps_2812 = A[12] & B[16]; 
assign ps_2811 = A[11] & B[17]; 
assign ps_2810 = A[10] & B[18]; 
assign ps_289 = A[9] & B[19]; 
assign ps_288 = A[8] & B[20]; 
assign ps_287 = A[7] & B[21]; 
assign ps_286 = A[6] & B[22]; 
assign ps_285 = A[5] & B[23]; 
assign ps_284 = A[4] & B[24]; 
assign ps_283 = A[3] & B[25]; 
assign ps_282 = A[2] & B[26]; 
assign ps_281 = A[1] & B[27]; 
assign ps_280 = A[0] & B[28]; 
assign ps_2929 = A[29] & B[0]; 
assign ps_2928 = A[28] & B[1]; 
assign ps_2927 = A[27] & B[2]; 
assign ps_2926 = A[26] & B[3]; 
assign ps_2925 = A[25] & B[4]; 
assign ps_2924 = A[24] & B[5]; 
assign ps_2923 = A[23] & B[6]; 
assign ps_2922 = A[22] & B[7]; 
assign ps_2921 = A[21] & B[8]; 
assign ps_2920 = A[20] & B[9]; 
assign ps_2919 = A[19] & B[10]; 
assign ps_2918 = A[18] & B[11]; 
assign ps_2917 = A[17] & B[12]; 
assign ps_2916 = A[16] & B[13]; 
assign ps_2915 = A[15] & B[14]; 
assign ps_2914 = A[14] & B[15]; 
assign ps_2913 = A[13] & B[16]; 
assign ps_2912 = A[12] & B[17]; 
assign ps_2911 = A[11] & B[18]; 
assign ps_2910 = A[10] & B[19]; 
assign ps_299 = A[9] & B[20]; 
assign ps_298 = A[8] & B[21]; 
assign ps_297 = A[7] & B[22]; 
assign ps_296 = A[6] & B[23]; 
assign ps_295 = A[5] & B[24]; 
assign ps_294 = A[4] & B[25]; 
assign ps_293 = A[3] & B[26]; 
assign ps_292 = A[2] & B[27]; 
assign ps_291 = A[1] & B[28]; 
assign ps_290 = A[0] & B[29]; 
assign ps_3030 = A[30] & B[0]; 
assign ps_3029 = A[29] & B[1]; 
assign ps_3028 = A[28] & B[2]; 
assign ps_3027 = A[27] & B[3]; 
assign ps_3026 = A[26] & B[4]; 
assign ps_3025 = A[25] & B[5]; 
assign ps_3024 = A[24] & B[6]; 
assign ps_3023 = A[23] & B[7]; 
assign ps_3022 = A[22] & B[8]; 
assign ps_3021 = A[21] & B[9]; 
assign ps_3020 = A[20] & B[10]; 
assign ps_3019 = A[19] & B[11]; 
assign ps_3018 = A[18] & B[12]; 
assign ps_3017 = A[17] & B[13]; 
assign ps_3016 = A[16] & B[14]; 
assign ps_3015 = A[15] & B[15]; 
assign ps_3014 = A[14] & B[16]; 
assign ps_3013 = A[13] & B[17]; 
assign ps_3012 = A[12] & B[18]; 
assign ps_3011 = A[11] & B[19]; 
assign ps_3010 = A[10] & B[20]; 
assign ps_309 = A[9] & B[21]; 
assign ps_308 = A[8] & B[22]; 
assign ps_307 = A[7] & B[23]; 
assign ps_306 = A[6] & B[24]; 
assign ps_305 = A[5] & B[25]; 
assign ps_304 = A[4] & B[26]; 
assign ps_303 = A[3] & B[27]; 
assign ps_302 = A[2] & B[28]; 
assign ps_301 = A[1] & B[29]; 
assign ps_300 = A[0] & B[30]; 
assign ps_3131 = A[31] & B[0]; 
assign ps_3130 = A[30] & B[1]; 
assign ps_3129 = A[29] & B[2]; 
assign ps_3128 = A[28] & B[3]; 
assign ps_3127 = A[27] & B[4]; 
assign ps_3126 = A[26] & B[5]; 
assign ps_3125 = A[25] & B[6]; 
assign ps_3124 = A[24] & B[7]; 
assign ps_3123 = A[23] & B[8]; 
assign ps_3122 = A[22] & B[9]; 
assign ps_3121 = A[21] & B[10]; 
assign ps_3120 = A[20] & B[11]; 
assign ps_3119 = A[19] & B[12]; 
assign ps_3118 = A[18] & B[13]; 
assign ps_3117 = A[17] & B[14]; 
assign ps_3116 = A[16] & B[15]; 
assign ps_3115 = A[15] & B[16]; 
assign ps_3114 = A[14] & B[17]; 
assign ps_3113 = A[13] & B[18]; 
assign ps_3112 = A[12] & B[19]; 
assign ps_3111 = A[11] & B[20]; 
assign ps_3110 = A[10] & B[21]; 
assign ps_319 = A[9] & B[22]; 
assign ps_318 = A[8] & B[23]; 
assign ps_317 = A[7] & B[24]; 
assign ps_316 = A[6] & B[25]; 
assign ps_315 = A[5] & B[26]; 
assign ps_314 = A[4] & B[27]; 
assign ps_313 = A[3] & B[28]; 
assign ps_312 = A[2] & B[29]; 
assign ps_311 = A[1] & B[30]; 
assign ps_310 = A[0] & B[31]; 
assign ps_3231 = A[31] & B[1]; 
assign ps_3230 = A[30] & B[2]; 
assign ps_3229 = A[29] & B[3]; 
assign ps_3228 = A[28] & B[4]; 
assign ps_3227 = A[27] & B[5]; 
assign ps_3226 = A[26] & B[6]; 
assign ps_3225 = A[25] & B[7]; 
assign ps_3224 = A[24] & B[8]; 
assign ps_3223 = A[23] & B[9]; 
assign ps_3222 = A[22] & B[10]; 
assign ps_3221 = A[21] & B[11]; 
assign ps_3220 = A[20] & B[12]; 
assign ps_3219 = A[19] & B[13]; 
assign ps_3218 = A[18] & B[14]; 
assign ps_3217 = A[17] & B[15]; 
assign ps_3216 = A[16] & B[16]; 
assign ps_3215 = A[15] & B[17]; 
assign ps_3214 = A[14] & B[18]; 
assign ps_3213 = A[13] & B[19]; 
assign ps_3212 = A[12] & B[20]; 
assign ps_3211 = A[11] & B[21]; 
assign ps_3210 = A[10] & B[22]; 
assign ps_329 = A[9] & B[23]; 
assign ps_328 = A[8] & B[24]; 
assign ps_327 = A[7] & B[25]; 
assign ps_326 = A[6] & B[26]; 
assign ps_325 = A[5] & B[27]; 
assign ps_324 = A[4] & B[28]; 
assign ps_323 = A[3] & B[29]; 
assign ps_322 = A[2] & B[30]; 
assign ps_321 = A[1] & B[31]; 
assign ps_3331 = A[31] & B[2]; 
assign ps_3330 = A[30] & B[3]; 
assign ps_3329 = A[29] & B[4]; 
assign ps_3328 = A[28] & B[5]; 
assign ps_3327 = A[27] & B[6]; 
assign ps_3326 = A[26] & B[7]; 
assign ps_3325 = A[25] & B[8]; 
assign ps_3324 = A[24] & B[9]; 
assign ps_3323 = A[23] & B[10]; 
assign ps_3322 = A[22] & B[11]; 
assign ps_3321 = A[21] & B[12]; 
assign ps_3320 = A[20] & B[13]; 
assign ps_3319 = A[19] & B[14]; 
assign ps_3318 = A[18] & B[15]; 
assign ps_3317 = A[17] & B[16]; 
assign ps_3316 = A[16] & B[17]; 
assign ps_3315 = A[15] & B[18]; 
assign ps_3314 = A[14] & B[19]; 
assign ps_3313 = A[13] & B[20]; 
assign ps_3312 = A[12] & B[21]; 
assign ps_3311 = A[11] & B[22]; 
assign ps_3310 = A[10] & B[23]; 
assign ps_339 = A[9] & B[24]; 
assign ps_338 = A[8] & B[25]; 
assign ps_337 = A[7] & B[26]; 
assign ps_336 = A[6] & B[27]; 
assign ps_335 = A[5] & B[28]; 
assign ps_334 = A[4] & B[29]; 
assign ps_333 = A[3] & B[30]; 
assign ps_332 = A[2] & B[31]; 
assign ps_3431 = A[31] & B[3]; 
assign ps_3430 = A[30] & B[4]; 
assign ps_3429 = A[29] & B[5]; 
assign ps_3428 = A[28] & B[6]; 
assign ps_3427 = A[27] & B[7]; 
assign ps_3426 = A[26] & B[8]; 
assign ps_3425 = A[25] & B[9]; 
assign ps_3424 = A[24] & B[10]; 
assign ps_3423 = A[23] & B[11]; 
assign ps_3422 = A[22] & B[12]; 
assign ps_3421 = A[21] & B[13]; 
assign ps_3420 = A[20] & B[14]; 
assign ps_3419 = A[19] & B[15]; 
assign ps_3418 = A[18] & B[16]; 
assign ps_3417 = A[17] & B[17]; 
assign ps_3416 = A[16] & B[18]; 
assign ps_3415 = A[15] & B[19]; 
assign ps_3414 = A[14] & B[20]; 
assign ps_3413 = A[13] & B[21]; 
assign ps_3412 = A[12] & B[22]; 
assign ps_3411 = A[11] & B[23]; 
assign ps_3410 = A[10] & B[24]; 
assign ps_349 = A[9] & B[25]; 
assign ps_348 = A[8] & B[26]; 
assign ps_347 = A[7] & B[27]; 
assign ps_346 = A[6] & B[28]; 
assign ps_345 = A[5] & B[29]; 
assign ps_344 = A[4] & B[30]; 
assign ps_343 = A[3] & B[31]; 
assign ps_3531 = A[31] & B[4]; 
assign ps_3530 = A[30] & B[5]; 
assign ps_3529 = A[29] & B[6]; 
assign ps_3528 = A[28] & B[7]; 
assign ps_3527 = A[27] & B[8]; 
assign ps_3526 = A[26] & B[9]; 
assign ps_3525 = A[25] & B[10]; 
assign ps_3524 = A[24] & B[11]; 
assign ps_3523 = A[23] & B[12]; 
assign ps_3522 = A[22] & B[13]; 
assign ps_3521 = A[21] & B[14]; 
assign ps_3520 = A[20] & B[15]; 
assign ps_3519 = A[19] & B[16]; 
assign ps_3518 = A[18] & B[17]; 
assign ps_3517 = A[17] & B[18]; 
assign ps_3516 = A[16] & B[19]; 
assign ps_3515 = A[15] & B[20]; 
assign ps_3514 = A[14] & B[21]; 
assign ps_3513 = A[13] & B[22]; 
assign ps_3512 = A[12] & B[23]; 
assign ps_3511 = A[11] & B[24]; 
assign ps_3510 = A[10] & B[25]; 
assign ps_359 = A[9] & B[26]; 
assign ps_358 = A[8] & B[27]; 
assign ps_357 = A[7] & B[28]; 
assign ps_356 = A[6] & B[29]; 
assign ps_355 = A[5] & B[30]; 
assign ps_354 = A[4] & B[31]; 
assign ps_3631 = A[31] & B[5]; 
assign ps_3630 = A[30] & B[6]; 
assign ps_3629 = A[29] & B[7]; 
assign ps_3628 = A[28] & B[8]; 
assign ps_3627 = A[27] & B[9]; 
assign ps_3626 = A[26] & B[10]; 
assign ps_3625 = A[25] & B[11]; 
assign ps_3624 = A[24] & B[12]; 
assign ps_3623 = A[23] & B[13]; 
assign ps_3622 = A[22] & B[14]; 
assign ps_3621 = A[21] & B[15]; 
assign ps_3620 = A[20] & B[16]; 
assign ps_3619 = A[19] & B[17]; 
assign ps_3618 = A[18] & B[18]; 
assign ps_3617 = A[17] & B[19]; 
assign ps_3616 = A[16] & B[20]; 
assign ps_3615 = A[15] & B[21]; 
assign ps_3614 = A[14] & B[22]; 
assign ps_3613 = A[13] & B[23]; 
assign ps_3612 = A[12] & B[24]; 
assign ps_3611 = A[11] & B[25]; 
assign ps_3610 = A[10] & B[26]; 
assign ps_369 = A[9] & B[27]; 
assign ps_368 = A[8] & B[28]; 
assign ps_367 = A[7] & B[29]; 
assign ps_366 = A[6] & B[30]; 
assign ps_365 = A[5] & B[31]; 
assign ps_3731 = A[31] & B[6]; 
assign ps_3730 = A[30] & B[7]; 
assign ps_3729 = A[29] & B[8]; 
assign ps_3728 = A[28] & B[9]; 
assign ps_3727 = A[27] & B[10]; 
assign ps_3726 = A[26] & B[11]; 
assign ps_3725 = A[25] & B[12]; 
assign ps_3724 = A[24] & B[13]; 
assign ps_3723 = A[23] & B[14]; 
assign ps_3722 = A[22] & B[15]; 
assign ps_3721 = A[21] & B[16]; 
assign ps_3720 = A[20] & B[17]; 
assign ps_3719 = A[19] & B[18]; 
assign ps_3718 = A[18] & B[19]; 
assign ps_3717 = A[17] & B[20]; 
assign ps_3716 = A[16] & B[21]; 
assign ps_3715 = A[15] & B[22]; 
assign ps_3714 = A[14] & B[23]; 
assign ps_3713 = A[13] & B[24]; 
assign ps_3712 = A[12] & B[25]; 
assign ps_3711 = A[11] & B[26]; 
assign ps_3710 = A[10] & B[27]; 
assign ps_379 = A[9] & B[28]; 
assign ps_378 = A[8] & B[29]; 
assign ps_377 = A[7] & B[30]; 
assign ps_376 = A[6] & B[31]; 
assign ps_3831 = A[31] & B[7]; 
assign ps_3830 = A[30] & B[8]; 
assign ps_3829 = A[29] & B[9]; 
assign ps_3828 = A[28] & B[10]; 
assign ps_3827 = A[27] & B[11]; 
assign ps_3826 = A[26] & B[12]; 
assign ps_3825 = A[25] & B[13]; 
assign ps_3824 = A[24] & B[14]; 
assign ps_3823 = A[23] & B[15]; 
assign ps_3822 = A[22] & B[16]; 
assign ps_3821 = A[21] & B[17]; 
assign ps_3820 = A[20] & B[18]; 
assign ps_3819 = A[19] & B[19]; 
assign ps_3818 = A[18] & B[20]; 
assign ps_3817 = A[17] & B[21]; 
assign ps_3816 = A[16] & B[22]; 
assign ps_3815 = A[15] & B[23]; 
assign ps_3814 = A[14] & B[24]; 
assign ps_3813 = A[13] & B[25]; 
assign ps_3812 = A[12] & B[26]; 
assign ps_3811 = A[11] & B[27]; 
assign ps_3810 = A[10] & B[28]; 
assign ps_389 = A[9] & B[29]; 
assign ps_388 = A[8] & B[30]; 
assign ps_387 = A[7] & B[31]; 
assign ps_3931 = A[31] & B[8]; 
assign ps_3930 = A[30] & B[9]; 
assign ps_3929 = A[29] & B[10]; 
assign ps_3928 = A[28] & B[11]; 
assign ps_3927 = A[27] & B[12]; 
assign ps_3926 = A[26] & B[13]; 
assign ps_3925 = A[25] & B[14]; 
assign ps_3924 = A[24] & B[15]; 
assign ps_3923 = A[23] & B[16]; 
assign ps_3922 = A[22] & B[17]; 
assign ps_3921 = A[21] & B[18]; 
assign ps_3920 = A[20] & B[19]; 
assign ps_3919 = A[19] & B[20]; 
assign ps_3918 = A[18] & B[21]; 
assign ps_3917 = A[17] & B[22]; 
assign ps_3916 = A[16] & B[23]; 
assign ps_3915 = A[15] & B[24]; 
assign ps_3914 = A[14] & B[25]; 
assign ps_3913 = A[13] & B[26]; 
assign ps_3912 = A[12] & B[27]; 
assign ps_3911 = A[11] & B[28]; 
assign ps_3910 = A[10] & B[29]; 
assign ps_399 = A[9] & B[30]; 
assign ps_398 = A[8] & B[31]; 
assign ps_4031 = A[31] & B[9]; 
assign ps_4030 = A[30] & B[10]; 
assign ps_4029 = A[29] & B[11]; 
assign ps_4028 = A[28] & B[12]; 
assign ps_4027 = A[27] & B[13]; 
assign ps_4026 = A[26] & B[14]; 
assign ps_4025 = A[25] & B[15]; 
assign ps_4024 = A[24] & B[16]; 
assign ps_4023 = A[23] & B[17]; 
assign ps_4022 = A[22] & B[18]; 
assign ps_4021 = A[21] & B[19]; 
assign ps_4020 = A[20] & B[20]; 
assign ps_4019 = A[19] & B[21]; 
assign ps_4018 = A[18] & B[22]; 
assign ps_4017 = A[17] & B[23]; 
assign ps_4016 = A[16] & B[24]; 
assign ps_4015 = A[15] & B[25]; 
assign ps_4014 = A[14] & B[26]; 
assign ps_4013 = A[13] & B[27]; 
assign ps_4012 = A[12] & B[28]; 
assign ps_4011 = A[11] & B[29]; 
assign ps_4010 = A[10] & B[30]; 
assign ps_409 = A[9] & B[31]; 
assign ps_4131 = A[31] & B[10]; 
assign ps_4130 = A[30] & B[11]; 
assign ps_4129 = A[29] & B[12]; 
assign ps_4128 = A[28] & B[13]; 
assign ps_4127 = A[27] & B[14]; 
assign ps_4126 = A[26] & B[15]; 
assign ps_4125 = A[25] & B[16]; 
assign ps_4124 = A[24] & B[17]; 
assign ps_4123 = A[23] & B[18]; 
assign ps_4122 = A[22] & B[19]; 
assign ps_4121 = A[21] & B[20]; 
assign ps_4120 = A[20] & B[21]; 
assign ps_4119 = A[19] & B[22]; 
assign ps_4118 = A[18] & B[23]; 
assign ps_4117 = A[17] & B[24]; 
assign ps_4116 = A[16] & B[25]; 
assign ps_4115 = A[15] & B[26]; 
assign ps_4114 = A[14] & B[27]; 
assign ps_4113 = A[13] & B[28]; 
assign ps_4112 = A[12] & B[29]; 
assign ps_4111 = A[11] & B[30]; 
assign ps_4110 = A[10] & B[31]; 
assign ps_4231 = A[31] & B[11]; 
assign ps_4230 = A[30] & B[12]; 
assign ps_4229 = A[29] & B[13]; 
assign ps_4228 = A[28] & B[14]; 
assign ps_4227 = A[27] & B[15]; 
assign ps_4226 = A[26] & B[16]; 
assign ps_4225 = A[25] & B[17]; 
assign ps_4224 = A[24] & B[18]; 
assign ps_4223 = A[23] & B[19]; 
assign ps_4222 = A[22] & B[20]; 
assign ps_4221 = A[21] & B[21]; 
assign ps_4220 = A[20] & B[22]; 
assign ps_4219 = A[19] & B[23]; 
assign ps_4218 = A[18] & B[24]; 
assign ps_4217 = A[17] & B[25]; 
assign ps_4216 = A[16] & B[26]; 
assign ps_4215 = A[15] & B[27]; 
assign ps_4214 = A[14] & B[28]; 
assign ps_4213 = A[13] & B[29]; 
assign ps_4212 = A[12] & B[30]; 
assign ps_4211 = A[11] & B[31]; 
assign ps_4331 = A[31] & B[12]; 
assign ps_4330 = A[30] & B[13]; 
assign ps_4329 = A[29] & B[14]; 
assign ps_4328 = A[28] & B[15]; 
assign ps_4327 = A[27] & B[16]; 
assign ps_4326 = A[26] & B[17]; 
assign ps_4325 = A[25] & B[18]; 
assign ps_4324 = A[24] & B[19]; 
assign ps_4323 = A[23] & B[20]; 
assign ps_4322 = A[22] & B[21]; 
assign ps_4321 = A[21] & B[22]; 
assign ps_4320 = A[20] & B[23]; 
assign ps_4319 = A[19] & B[24]; 
assign ps_4318 = A[18] & B[25]; 
assign ps_4317 = A[17] & B[26]; 
assign ps_4316 = A[16] & B[27]; 
assign ps_4315 = A[15] & B[28]; 
assign ps_4314 = A[14] & B[29]; 
assign ps_4313 = A[13] & B[30]; 
assign ps_4312 = A[12] & B[31]; 
assign ps_4431 = A[31] & B[13]; 
assign ps_4430 = A[30] & B[14]; 
assign ps_4429 = A[29] & B[15]; 
assign ps_4428 = A[28] & B[16]; 
assign ps_4427 = A[27] & B[17]; 
assign ps_4426 = A[26] & B[18]; 
assign ps_4425 = A[25] & B[19]; 
assign ps_4424 = A[24] & B[20]; 
assign ps_4423 = A[23] & B[21]; 
assign ps_4422 = A[22] & B[22]; 
assign ps_4421 = A[21] & B[23]; 
assign ps_4420 = A[20] & B[24]; 
assign ps_4419 = A[19] & B[25]; 
assign ps_4418 = A[18] & B[26]; 
assign ps_4417 = A[17] & B[27]; 
assign ps_4416 = A[16] & B[28]; 
assign ps_4415 = A[15] & B[29]; 
assign ps_4414 = A[14] & B[30]; 
assign ps_4413 = A[13] & B[31]; 
assign ps_4531 = A[31] & B[14]; 
assign ps_4530 = A[30] & B[15]; 
assign ps_4529 = A[29] & B[16]; 
assign ps_4528 = A[28] & B[17]; 
assign ps_4527 = A[27] & B[18]; 
assign ps_4526 = A[26] & B[19]; 
assign ps_4525 = A[25] & B[20]; 
assign ps_4524 = A[24] & B[21]; 
assign ps_4523 = A[23] & B[22]; 
assign ps_4522 = A[22] & B[23]; 
assign ps_4521 = A[21] & B[24]; 
assign ps_4520 = A[20] & B[25]; 
assign ps_4519 = A[19] & B[26]; 
assign ps_4518 = A[18] & B[27]; 
assign ps_4517 = A[17] & B[28]; 
assign ps_4516 = A[16] & B[29]; 
assign ps_4515 = A[15] & B[30]; 
assign ps_4514 = A[14] & B[31]; 
assign ps_4631 = A[31] & B[15]; 
assign ps_4630 = A[30] & B[16]; 
assign ps_4629 = A[29] & B[17]; 
assign ps_4628 = A[28] & B[18]; 
assign ps_4627 = A[27] & B[19]; 
assign ps_4626 = A[26] & B[20]; 
assign ps_4625 = A[25] & B[21]; 
assign ps_4624 = A[24] & B[22]; 
assign ps_4623 = A[23] & B[23]; 
assign ps_4622 = A[22] & B[24]; 
assign ps_4621 = A[21] & B[25]; 
assign ps_4620 = A[20] & B[26]; 
assign ps_4619 = A[19] & B[27]; 
assign ps_4618 = A[18] & B[28]; 
assign ps_4617 = A[17] & B[29]; 
assign ps_4616 = A[16] & B[30]; 
assign ps_4615 = A[15] & B[31]; 
assign ps_4731 = A[31] & B[16]; 
assign ps_4730 = A[30] & B[17]; 
assign ps_4729 = A[29] & B[18]; 
assign ps_4728 = A[28] & B[19]; 
assign ps_4727 = A[27] & B[20]; 
assign ps_4726 = A[26] & B[21]; 
assign ps_4725 = A[25] & B[22]; 
assign ps_4724 = A[24] & B[23]; 
assign ps_4723 = A[23] & B[24]; 
assign ps_4722 = A[22] & B[25]; 
assign ps_4721 = A[21] & B[26]; 
assign ps_4720 = A[20] & B[27]; 
assign ps_4719 = A[19] & B[28]; 
assign ps_4718 = A[18] & B[29]; 
assign ps_4717 = A[17] & B[30]; 
assign ps_4716 = A[16] & B[31]; 
assign ps_4831 = A[31] & B[17]; 
assign ps_4830 = A[30] & B[18]; 
assign ps_4829 = A[29] & B[19]; 
assign ps_4828 = A[28] & B[20]; 
assign ps_4827 = A[27] & B[21]; 
assign ps_4826 = A[26] & B[22]; 
assign ps_4825 = A[25] & B[23]; 
assign ps_4824 = A[24] & B[24]; 
assign ps_4823 = A[23] & B[25]; 
assign ps_4822 = A[22] & B[26]; 
assign ps_4821 = A[21] & B[27]; 
assign ps_4820 = A[20] & B[28]; 
assign ps_4819 = A[19] & B[29]; 
assign ps_4818 = A[18] & B[30]; 
assign ps_4817 = A[17] & B[31]; 
assign ps_4931 = A[31] & B[18]; 
assign ps_4930 = A[30] & B[19]; 
assign ps_4929 = A[29] & B[20]; 
assign ps_4928 = A[28] & B[21]; 
assign ps_4927 = A[27] & B[22]; 
assign ps_4926 = A[26] & B[23]; 
assign ps_4925 = A[25] & B[24]; 
assign ps_4924 = A[24] & B[25]; 
assign ps_4923 = A[23] & B[26]; 
assign ps_4922 = A[22] & B[27]; 
assign ps_4921 = A[21] & B[28]; 
assign ps_4920 = A[20] & B[29]; 
assign ps_4919 = A[19] & B[30]; 
assign ps_4918 = A[18] & B[31]; 
assign ps_5031 = A[31] & B[19]; 
assign ps_5030 = A[30] & B[20]; 
assign ps_5029 = A[29] & B[21]; 
assign ps_5028 = A[28] & B[22]; 
assign ps_5027 = A[27] & B[23]; 
assign ps_5026 = A[26] & B[24]; 
assign ps_5025 = A[25] & B[25]; 
assign ps_5024 = A[24] & B[26]; 
assign ps_5023 = A[23] & B[27]; 
assign ps_5022 = A[22] & B[28]; 
assign ps_5021 = A[21] & B[29]; 
assign ps_5020 = A[20] & B[30]; 
assign ps_5019 = A[19] & B[31]; 
assign ps_5131 = A[31] & B[20]; 
assign ps_5130 = A[30] & B[21]; 
assign ps_5129 = A[29] & B[22]; 
assign ps_5128 = A[28] & B[23]; 
assign ps_5127 = A[27] & B[24]; 
assign ps_5126 = A[26] & B[25]; 
assign ps_5125 = A[25] & B[26]; 
assign ps_5124 = A[24] & B[27]; 
assign ps_5123 = A[23] & B[28]; 
assign ps_5122 = A[22] & B[29]; 
assign ps_5121 = A[21] & B[30]; 
assign ps_5120 = A[20] & B[31]; 
assign ps_5231 = A[31] & B[21]; 
assign ps_5230 = A[30] & B[22]; 
assign ps_5229 = A[29] & B[23]; 
assign ps_5228 = A[28] & B[24]; 
assign ps_5227 = A[27] & B[25]; 
assign ps_5226 = A[26] & B[26]; 
assign ps_5225 = A[25] & B[27]; 
assign ps_5224 = A[24] & B[28]; 
assign ps_5223 = A[23] & B[29]; 
assign ps_5222 = A[22] & B[30]; 
assign ps_5221 = A[21] & B[31]; 
assign ps_5331 = A[31] & B[22]; 
assign ps_5330 = A[30] & B[23]; 
assign ps_5329 = A[29] & B[24]; 
assign ps_5328 = A[28] & B[25]; 
assign ps_5327 = A[27] & B[26]; 
assign ps_5326 = A[26] & B[27]; 
assign ps_5325 = A[25] & B[28]; 
assign ps_5324 = A[24] & B[29]; 
assign ps_5323 = A[23] & B[30]; 
assign ps_5322 = A[22] & B[31]; 
assign ps_5431 = A[31] & B[23]; 
assign ps_5430 = A[30] & B[24]; 
assign ps_5429 = A[29] & B[25]; 
assign ps_5428 = A[28] & B[26]; 
assign ps_5427 = A[27] & B[27]; 
assign ps_5426 = A[26] & B[28]; 
assign ps_5425 = A[25] & B[29]; 
assign ps_5424 = A[24] & B[30]; 
assign ps_5423 = A[23] & B[31]; 
assign ps_5531 = A[31] & B[24]; 
assign ps_5530 = A[30] & B[25]; 
assign ps_5529 = A[29] & B[26]; 
assign ps_5528 = A[28] & B[27]; 
assign ps_5527 = A[27] & B[28]; 
assign ps_5526 = A[26] & B[29]; 
assign ps_5525 = A[25] & B[30]; 
assign ps_5524 = A[24] & B[31]; 
assign ps_5631 = A[31] & B[25]; 
assign ps_5630 = A[30] & B[26]; 
assign ps_5629 = A[29] & B[27]; 
assign ps_5628 = A[28] & B[28]; 
assign ps_5627 = A[27] & B[29]; 
assign ps_5626 = A[26] & B[30]; 
assign ps_5625 = A[25] & B[31]; 
assign ps_5731 = A[31] & B[26]; 
assign ps_5730 = A[30] & B[27]; 
assign ps_5729 = A[29] & B[28]; 
assign ps_5728 = A[28] & B[29]; 
assign ps_5727 = A[27] & B[30]; 
assign ps_5726 = A[26] & B[31]; 
assign ps_5831 = A[31] & B[27]; 
assign ps_5830 = A[30] & B[28]; 
assign ps_5829 = A[29] & B[29]; 
assign ps_5828 = A[28] & B[30]; 
assign ps_5827 = A[27] & B[31]; 
assign ps_5931 = A[31] & B[28]; 
assign ps_5930 = A[30] & B[29]; 
assign ps_5929 = A[29] & B[30]; 
assign ps_5928 = A[28] & B[31]; 
assign ps_6031 = A[31] & B[29]; 
assign ps_6030 = A[30] & B[30]; 
assign ps_6029 = A[29] & B[31]; 
assign ps_6131 = A[31] & B[30]; 
assign ps_6130 = A[30] & B[31]; 
assign ps_6231 = A[31] & B[31]; 
logic s1_280_hacout, s1_280_has, s1_290_facout, s1_290_fas, s1_290_hacout, s1_290_has, s1_300_facout, s1_300_fas, s1_301_facout, s1_301_fas, s1_300_hacout, s1_300_has, s1_310_facout, s1_310_fas, s1_311_facout, s1_311_fas, s1_312_facout, s1_312_fas, s1_310_hacout, s1_310_has, s1_320_facout, s1_320_fas, s1_321_facout, s1_321_fas, s1_322_facout, s1_322_fas, s1_320_hacout, s1_320_has, s1_330_facout, s1_330_fas, s1_331_facout, s1_331_fas, s1_332_facout, s1_332_fas, s1_340_facout, s1_340_fas, s1_341_facout, s1_341_fas, s1_350_facout, s1_350_fas;
/* ========================= Stage 1 ========================= */
half_adder s1_28ha0 ( .A(ps_2828), .B(ps_2827), .S(s1_280_has), .Cout(s1_280_hacout));
full_adder s1_29fa0 ( .A(ps_2929), .B(ps_2928), .Cin(ps_2927), .S(s1_290_fas), .Cout(s1_290_facout));
half_adder s1_29ha0 ( .A(ps_2926), .B(ps_2925), .S(s1_290_has), .Cout(s1_290_hacout));
full_adder s1_30fa0 ( .A(ps_3030), .B(ps_3029), .Cin(ps_3028), .S(s1_300_fas), .Cout(s1_300_facout));
full_adder s1_30fa1 ( .A(ps_3027), .B(ps_3026), .Cin(ps_3025), .S(s1_301_fas), .Cout(s1_301_facout));
half_adder s1_30ha0 ( .A(ps_3024), .B(ps_3023), .S(s1_300_has), .Cout(s1_300_hacout));
full_adder s1_31fa0 ( .A(ps_3131), .B(ps_3130), .Cin(ps_3129), .S(s1_310_fas), .Cout(s1_310_facout));
full_adder s1_31fa1 ( .A(ps_3128), .B(ps_3127), .Cin(ps_3126), .S(s1_311_fas), .Cout(s1_311_facout));
full_adder s1_31fa2 ( .A(ps_3125), .B(ps_3124), .Cin(ps_3123), .S(s1_312_fas), .Cout(s1_312_facout));
half_adder s1_31ha0 ( .A(ps_3122), .B(ps_3121), .S(s1_310_has), .Cout(s1_310_hacout));
full_adder s1_32fa0 ( .A(ps_3231), .B(ps_3230), .Cin(ps_3229), .S(s1_320_fas), .Cout(s1_320_facout));
full_adder s1_32fa1 ( .A(ps_3228), .B(ps_3227), .Cin(ps_3226), .S(s1_321_fas), .Cout(s1_321_facout));
full_adder s1_32fa2 ( .A(ps_3225), .B(ps_3224), .Cin(ps_3223), .S(s1_322_fas), .Cout(s1_322_facout));
half_adder s1_32ha0 ( .A(ps_3222), .B(ps_3221), .S(s1_320_has), .Cout(s1_320_hacout));
full_adder s1_33fa0 ( .A(ps_3331), .B(ps_3330), .Cin(ps_3329), .S(s1_330_fas), .Cout(s1_330_facout));
full_adder s1_33fa1 ( .A(ps_3328), .B(ps_3327), .Cin(ps_3326), .S(s1_331_fas), .Cout(s1_331_facout));
full_adder s1_33fa2 ( .A(ps_3325), .B(ps_3324), .Cin(ps_3323), .S(s1_332_fas), .Cout(s1_332_facout));
full_adder s1_34fa0 ( .A(ps_3431), .B(ps_3430), .Cin(ps_3429), .S(s1_340_fas), .Cout(s1_340_facout));
full_adder s1_34fa1 ( .A(ps_3428), .B(ps_3427), .Cin(ps_3426), .S(s1_341_fas), .Cout(s1_341_facout));
full_adder s1_35fa0 ( .A(ps_3531), .B(ps_3530), .Cin(ps_3529), .S(s1_350_fas), .Cout(s1_350_facout));
logic s2_190_hacout, s2_190_has, s2_200_facout, s2_200_fas, s2_200_hacout, s2_200_has, s2_210_facout, s2_210_fas, s2_211_facout, s2_211_fas, s2_210_hacout, s2_210_has, s2_220_facout, s2_220_fas, s2_221_facout, s2_221_fas, s2_222_facout, s2_222_fas, s2_220_hacout, s2_220_has, s2_230_facout, s2_230_fas, s2_231_facout, s2_231_fas, s2_232_facout, s2_232_fas, s2_233_facout, s2_233_fas, s2_230_hacout, s2_230_has, s2_240_facout, s2_240_fas, s2_241_facout, s2_241_fas, s2_242_facout, s2_242_fas, s2_243_facout, s2_243_fas, s2_244_facout, s2_244_fas, s2_240_hacout, s2_240_has, s2_250_facout, s2_250_fas, s2_251_facout, s2_251_fas, s2_252_facout, s2_252_fas, s2_253_facout, s2_253_fas, s2_254_facout, s2_254_fas, s2_255_facout, s2_255_fas, s2_250_hacout, s2_250_has, s2_260_facout, s2_260_fas, s2_261_facout, s2_261_fas, s2_262_facout, s2_262_fas, s2_263_facout, s2_263_fas, s2_264_facout, s2_264_fas, s2_265_facout, s2_265_fas, s2_266_facout, s2_266_fas, s2_260_hacout, s2_260_has, s2_270_facout, s2_270_fas, s2_271_facout, s2_271_fas, s2_272_facout, s2_272_fas, s2_273_facout, s2_273_fas, s2_274_facout, s2_274_fas, s2_275_facout, s2_275_fas, s2_276_facout, s2_276_fas, s2_277_facout, s2_277_fas, s2_270_hacout, s2_270_has, s2_280_facout, s2_280_fas, s2_281_facout, s2_281_fas, s2_282_facout, s2_282_fas, s2_283_facout, s2_283_fas, s2_284_facout, s2_284_fas, s2_285_facout, s2_285_fas, s2_286_facout, s2_286_fas, s2_287_facout, s2_287_fas, s2_288_facout, s2_288_fas, s2_290_facout, s2_290_fas, s2_291_facout, s2_291_fas, s2_292_facout, s2_292_fas, s2_293_facout, s2_293_fas, s2_294_facout, s2_294_fas, s2_295_facout, s2_295_fas, s2_296_facout, s2_296_fas, s2_297_facout, s2_297_fas, s2_298_facout, s2_298_fas, s2_300_facout, s2_300_fas, s2_301_facout, s2_301_fas, s2_302_facout, s2_302_fas, s2_303_facout, s2_303_fas, s2_304_facout, s2_304_fas, s2_305_facout, s2_305_fas, s2_306_facout, s2_306_fas, s2_307_facout, s2_307_fas, s2_308_facout, s2_308_fas, s2_310_facout, s2_310_fas, s2_311_facout, s2_311_fas, s2_312_facout, s2_312_fas, s2_313_facout, s2_313_fas, s2_314_facout, s2_314_fas, s2_315_facout, s2_315_fas, s2_316_facout, s2_316_fas, s2_317_facout, s2_317_fas, s2_318_facout, s2_318_fas, s2_320_facout, s2_320_fas, s2_321_facout, s2_321_fas, s2_322_facout, s2_322_fas, s2_323_facout, s2_323_fas, s2_324_facout, s2_324_fas, s2_325_facout, s2_325_fas, s2_326_facout, s2_326_fas, s2_327_facout, s2_327_fas, s2_328_facout, s2_328_fas, s2_330_facout, s2_330_fas, s2_331_facout, s2_331_fas, s2_332_facout, s2_332_fas, s2_333_facout, s2_333_fas, s2_334_facout, s2_334_fas, s2_335_facout, s2_335_fas, s2_336_facout, s2_336_fas, s2_337_facout, s2_337_fas, s2_338_facout, s2_338_fas, s2_340_facout, s2_340_fas, s2_341_facout, s2_341_fas, s2_342_facout, s2_342_fas, s2_343_facout, s2_343_fas, s2_344_facout, s2_344_fas, s2_345_facout, s2_345_fas, s2_346_facout, s2_346_fas, s2_347_facout, s2_347_fas, s2_348_facout, s2_348_fas, s2_350_facout, s2_350_fas, s2_351_facout, s2_351_fas, s2_352_facout, s2_352_fas, s2_353_facout, s2_353_fas, s2_354_facout, s2_354_fas, s2_355_facout, s2_355_fas, s2_356_facout, s2_356_fas, s2_357_facout, s2_357_fas, s2_358_facout, s2_358_fas, s2_360_facout, s2_360_fas, s2_361_facout, s2_361_fas, s2_362_facout, s2_362_fas, s2_363_facout, s2_363_fas, s2_364_facout, s2_364_fas, s2_365_facout, s2_365_fas, s2_366_facout, s2_366_fas, s2_367_facout, s2_367_fas, s2_368_facout, s2_368_fas, s2_370_facout, s2_370_fas, s2_371_facout, s2_371_fas, s2_372_facout, s2_372_fas, s2_373_facout, s2_373_fas, s2_374_facout, s2_374_fas, s2_375_facout, s2_375_fas, s2_376_facout, s2_376_fas, s2_377_facout, s2_377_fas, s2_380_facout, s2_380_fas, s2_381_facout, s2_381_fas, s2_382_facout, s2_382_fas, s2_383_facout, s2_383_fas, s2_384_facout, s2_384_fas, s2_385_facout, s2_385_fas, s2_386_facout, s2_386_fas, s2_390_facout, s2_390_fas, s2_391_facout, s2_391_fas, s2_392_facout, s2_392_fas, s2_393_facout, s2_393_fas, s2_394_facout, s2_394_fas, s2_395_facout, s2_395_fas, s2_400_facout, s2_400_fas, s2_401_facout, s2_401_fas, s2_402_facout, s2_402_fas, s2_403_facout, s2_403_fas, s2_404_facout, s2_404_fas, s2_410_facout, s2_410_fas, s2_411_facout, s2_411_fas, s2_412_facout, s2_412_fas, s2_413_facout, s2_413_fas, s2_420_facout, s2_420_fas, s2_421_facout, s2_421_fas, s2_422_facout, s2_422_fas, s2_430_facout, s2_430_fas, s2_431_facout, s2_431_fas, s2_440_facout, s2_440_fas;
/* ========================= Stage 2 ========================= */
half_adder s2_19ha0 ( .A(ps_1919), .B(ps_1918), .S(s2_190_has), .Cout(s2_190_hacout));
full_adder s2_20fa0 ( .A(ps_2020), .B(ps_2019), .Cin(ps_2018), .S(s2_200_fas), .Cout(s2_200_facout));
half_adder s2_20ha0 ( .A(ps_2017), .B(ps_2016), .S(s2_200_has), .Cout(s2_200_hacout));
full_adder s2_21fa0 ( .A(ps_2121), .B(ps_2120), .Cin(ps_2119), .S(s2_210_fas), .Cout(s2_210_facout));
full_adder s2_21fa1 ( .A(ps_2118), .B(ps_2117), .Cin(ps_2116), .S(s2_211_fas), .Cout(s2_211_facout));
half_adder s2_21ha0 ( .A(ps_2115), .B(ps_2114), .S(s2_210_has), .Cout(s2_210_hacout));
full_adder s2_22fa0 ( .A(ps_2222), .B(ps_2221), .Cin(ps_2220), .S(s2_220_fas), .Cout(s2_220_facout));
full_adder s2_22fa1 ( .A(ps_2219), .B(ps_2218), .Cin(ps_2217), .S(s2_221_fas), .Cout(s2_221_facout));
full_adder s2_22fa2 ( .A(ps_2216), .B(ps_2215), .Cin(ps_2214), .S(s2_222_fas), .Cout(s2_222_facout));
half_adder s2_22ha0 ( .A(ps_2213), .B(ps_2212), .S(s2_220_has), .Cout(s2_220_hacout));
full_adder s2_23fa0 ( .A(ps_2323), .B(ps_2322), .Cin(ps_2321), .S(s2_230_fas), .Cout(s2_230_facout));
full_adder s2_23fa1 ( .A(ps_2320), .B(ps_2319), .Cin(ps_2318), .S(s2_231_fas), .Cout(s2_231_facout));
full_adder s2_23fa2 ( .A(ps_2317), .B(ps_2316), .Cin(ps_2315), .S(s2_232_fas), .Cout(s2_232_facout));
full_adder s2_23fa3 ( .A(ps_2314), .B(ps_2313), .Cin(ps_2312), .S(s2_233_fas), .Cout(s2_233_facout));
half_adder s2_23ha0 ( .A(ps_2311), .B(ps_2310), .S(s2_230_has), .Cout(s2_230_hacout));
full_adder s2_24fa0 ( .A(ps_2424), .B(ps_2423), .Cin(ps_2422), .S(s2_240_fas), .Cout(s2_240_facout));
full_adder s2_24fa1 ( .A(ps_2421), .B(ps_2420), .Cin(ps_2419), .S(s2_241_fas), .Cout(s2_241_facout));
full_adder s2_24fa2 ( .A(ps_2418), .B(ps_2417), .Cin(ps_2416), .S(s2_242_fas), .Cout(s2_242_facout));
full_adder s2_24fa3 ( .A(ps_2415), .B(ps_2414), .Cin(ps_2413), .S(s2_243_fas), .Cout(s2_243_facout));
full_adder s2_24fa4 ( .A(ps_2412), .B(ps_2411), .Cin(ps_2410), .S(s2_244_fas), .Cout(s2_244_facout));
half_adder s2_24ha0 ( .A(ps_249), .B(ps_248), .S(s2_240_has), .Cout(s2_240_hacout));
full_adder s2_25fa0 ( .A(ps_2525), .B(ps_2524), .Cin(ps_2523), .S(s2_250_fas), .Cout(s2_250_facout));
full_adder s2_25fa1 ( .A(ps_2522), .B(ps_2521), .Cin(ps_2520), .S(s2_251_fas), .Cout(s2_251_facout));
full_adder s2_25fa2 ( .A(ps_2519), .B(ps_2518), .Cin(ps_2517), .S(s2_252_fas), .Cout(s2_252_facout));
full_adder s2_25fa3 ( .A(ps_2516), .B(ps_2515), .Cin(ps_2514), .S(s2_253_fas), .Cout(s2_253_facout));
full_adder s2_25fa4 ( .A(ps_2513), .B(ps_2512), .Cin(ps_2511), .S(s2_254_fas), .Cout(s2_254_facout));
full_adder s2_25fa5 ( .A(ps_2510), .B(ps_259), .Cin(ps_258), .S(s2_255_fas), .Cout(s2_255_facout));
half_adder s2_25ha0 ( .A(ps_257), .B(ps_256), .S(s2_250_has), .Cout(s2_250_hacout));
full_adder s2_26fa0 ( .A(ps_2626), .B(ps_2625), .Cin(ps_2624), .S(s2_260_fas), .Cout(s2_260_facout));
full_adder s2_26fa1 ( .A(ps_2623), .B(ps_2622), .Cin(ps_2621), .S(s2_261_fas), .Cout(s2_261_facout));
full_adder s2_26fa2 ( .A(ps_2620), .B(ps_2619), .Cin(ps_2618), .S(s2_262_fas), .Cout(s2_262_facout));
full_adder s2_26fa3 ( .A(ps_2617), .B(ps_2616), .Cin(ps_2615), .S(s2_263_fas), .Cout(s2_263_facout));
full_adder s2_26fa4 ( .A(ps_2614), .B(ps_2613), .Cin(ps_2612), .S(s2_264_fas), .Cout(s2_264_facout));
full_adder s2_26fa5 ( .A(ps_2611), .B(ps_2610), .Cin(ps_269), .S(s2_265_fas), .Cout(s2_265_facout));
full_adder s2_26fa6 ( .A(ps_268), .B(ps_267), .Cin(ps_266), .S(s2_266_fas), .Cout(s2_266_facout));
half_adder s2_26ha0 ( .A(ps_265), .B(ps_264), .S(s2_260_has), .Cout(s2_260_hacout));
full_adder s2_27fa0 ( .A(ps_2727), .B(ps_2726), .Cin(ps_2725), .S(s2_270_fas), .Cout(s2_270_facout));
full_adder s2_27fa1 ( .A(ps_2724), .B(ps_2723), .Cin(ps_2722), .S(s2_271_fas), .Cout(s2_271_facout));
full_adder s2_27fa2 ( .A(ps_2721), .B(ps_2720), .Cin(ps_2719), .S(s2_272_fas), .Cout(s2_272_facout));
full_adder s2_27fa3 ( .A(ps_2718), .B(ps_2717), .Cin(ps_2716), .S(s2_273_fas), .Cout(s2_273_facout));
full_adder s2_27fa4 ( .A(ps_2715), .B(ps_2714), .Cin(ps_2713), .S(s2_274_fas), .Cout(s2_274_facout));
full_adder s2_27fa5 ( .A(ps_2712), .B(ps_2711), .Cin(ps_2710), .S(s2_275_fas), .Cout(s2_275_facout));
full_adder s2_27fa6 ( .A(ps_279), .B(ps_278), .Cin(ps_277), .S(s2_276_fas), .Cout(s2_276_facout));
full_adder s2_27fa7 ( .A(ps_276), .B(ps_275), .Cin(ps_274), .S(s2_277_fas), .Cout(s2_277_facout));
half_adder s2_27ha0 ( .A(ps_273), .B(ps_272), .S(s2_270_has), .Cout(s2_270_hacout));
full_adder s2_28fa0 ( .A(ps_2826), .B(ps_2825), .Cin(ps_2824), .S(s2_280_fas), .Cout(s2_280_facout));
full_adder s2_28fa1 ( .A(ps_2823), .B(ps_2822), .Cin(ps_2821), .S(s2_281_fas), .Cout(s2_281_facout));
full_adder s2_28fa2 ( .A(ps_2820), .B(ps_2819), .Cin(ps_2818), .S(s2_282_fas), .Cout(s2_282_facout));
full_adder s2_28fa3 ( .A(ps_2817), .B(ps_2816), .Cin(ps_2815), .S(s2_283_fas), .Cout(s2_283_facout));
full_adder s2_28fa4 ( .A(ps_2814), .B(ps_2813), .Cin(ps_2812), .S(s2_284_fas), .Cout(s2_284_facout));
full_adder s2_28fa5 ( .A(ps_2811), .B(ps_2810), .Cin(ps_289), .S(s2_285_fas), .Cout(s2_285_facout));
full_adder s2_28fa6 ( .A(ps_288), .B(ps_287), .Cin(ps_286), .S(s2_286_fas), .Cout(s2_286_facout));
full_adder s2_28fa7 ( .A(ps_285), .B(ps_284), .Cin(ps_283), .S(s2_287_fas), .Cout(s2_287_facout));
full_adder s2_28fa8 ( .A(ps_282), .B(ps_281), .Cin(ps_280), .S(s2_288_fas), .Cout(s2_288_facout));
full_adder s2_29fa0 ( .A(ps_2924), .B(ps_2923), .Cin(ps_2922), .S(s2_290_fas), .Cout(s2_290_facout));
full_adder s2_29fa1 ( .A(ps_2921), .B(ps_2920), .Cin(ps_2919), .S(s2_291_fas), .Cout(s2_291_facout));
full_adder s2_29fa2 ( .A(ps_2918), .B(ps_2917), .Cin(ps_2916), .S(s2_292_fas), .Cout(s2_292_facout));
full_adder s2_29fa3 ( .A(ps_2915), .B(ps_2914), .Cin(ps_2913), .S(s2_293_fas), .Cout(s2_293_facout));
full_adder s2_29fa4 ( .A(ps_2912), .B(ps_2911), .Cin(ps_2910), .S(s2_294_fas), .Cout(s2_294_facout));
full_adder s2_29fa5 ( .A(ps_299), .B(ps_298), .Cin(ps_297), .S(s2_295_fas), .Cout(s2_295_facout));
full_adder s2_29fa6 ( .A(ps_296), .B(ps_295), .Cin(ps_294), .S(s2_296_fas), .Cout(s2_296_facout));
full_adder s2_29fa7 ( .A(ps_293), .B(ps_292), .Cin(ps_291), .S(s2_297_fas), .Cout(s2_297_facout));
full_adder s2_29fa8 ( .A(ps_290), .B(s1_280_hacout), .Cin(s1_290_fas), .S(s2_298_fas), .Cout(s2_298_facout));
full_adder s2_30fa0 ( .A(ps_3022), .B(ps_3021), .Cin(ps_3020), .S(s2_300_fas), .Cout(s2_300_facout));
full_adder s2_30fa1 ( .A(ps_3019), .B(ps_3018), .Cin(ps_3017), .S(s2_301_fas), .Cout(s2_301_facout));
full_adder s2_30fa2 ( .A(ps_3016), .B(ps_3015), .Cin(ps_3014), .S(s2_302_fas), .Cout(s2_302_facout));
full_adder s2_30fa3 ( .A(ps_3013), .B(ps_3012), .Cin(ps_3011), .S(s2_303_fas), .Cout(s2_303_facout));
full_adder s2_30fa4 ( .A(ps_3010), .B(ps_309), .Cin(ps_308), .S(s2_304_fas), .Cout(s2_304_facout));
full_adder s2_30fa5 ( .A(ps_307), .B(ps_306), .Cin(ps_305), .S(s2_305_fas), .Cout(s2_305_facout));
full_adder s2_30fa6 ( .A(ps_304), .B(ps_303), .Cin(ps_302), .S(s2_306_fas), .Cout(s2_306_facout));
full_adder s2_30fa7 ( .A(ps_301), .B(ps_300), .Cin(s1_290_facout), .S(s2_307_fas), .Cout(s2_307_facout));
full_adder s2_30fa8 ( .A(s1_290_hacout), .B(s1_300_fas), .Cin(s1_301_fas), .S(s2_308_fas), .Cout(s2_308_facout));
full_adder s2_31fa0 ( .A(ps_3120), .B(ps_3119), .Cin(ps_3118), .S(s2_310_fas), .Cout(s2_310_facout));
full_adder s2_31fa1 ( .A(ps_3117), .B(ps_3116), .Cin(ps_3115), .S(s2_311_fas), .Cout(s2_311_facout));
full_adder s2_31fa2 ( .A(ps_3114), .B(ps_3113), .Cin(ps_3112), .S(s2_312_fas), .Cout(s2_312_facout));
full_adder s2_31fa3 ( .A(ps_3111), .B(ps_3110), .Cin(ps_319), .S(s2_313_fas), .Cout(s2_313_facout));
full_adder s2_31fa4 ( .A(ps_318), .B(ps_317), .Cin(ps_316), .S(s2_314_fas), .Cout(s2_314_facout));
full_adder s2_31fa5 ( .A(ps_315), .B(ps_314), .Cin(ps_313), .S(s2_315_fas), .Cout(s2_315_facout));
full_adder s2_31fa6 ( .A(ps_312), .B(ps_311), .Cin(ps_310), .S(s2_316_fas), .Cout(s2_316_facout));
full_adder s2_31fa7 ( .A(s1_300_facout), .B(s1_301_facout), .Cin(s1_300_hacout), .S(s2_317_fas), .Cout(s2_317_facout));
full_adder s2_31fa8 ( .A(s1_310_fas), .B(s1_311_fas), .Cin(s1_312_fas), .S(s2_318_fas), .Cout(s2_318_facout));
full_adder s2_32fa0 ( .A(ps_3220), .B(ps_3219), .Cin(ps_3218), .S(s2_320_fas), .Cout(s2_320_facout));
full_adder s2_32fa1 ( .A(ps_3217), .B(ps_3216), .Cin(ps_3215), .S(s2_321_fas), .Cout(s2_321_facout));
full_adder s2_32fa2 ( .A(ps_3214), .B(ps_3213), .Cin(ps_3212), .S(s2_322_fas), .Cout(s2_322_facout));
full_adder s2_32fa3 ( .A(ps_3211), .B(ps_3210), .Cin(ps_329), .S(s2_323_fas), .Cout(s2_323_facout));
full_adder s2_32fa4 ( .A(ps_328), .B(ps_327), .Cin(ps_326), .S(s2_324_fas), .Cout(s2_324_facout));
full_adder s2_32fa5 ( .A(ps_325), .B(ps_324), .Cin(ps_323), .S(s2_325_fas), .Cout(s2_325_facout));
full_adder s2_32fa6 ( .A(ps_322), .B(ps_321), .Cin(s1_310_facout), .S(s2_326_fas), .Cout(s2_326_facout));
full_adder s2_32fa7 ( .A(s1_311_facout), .B(s1_312_facout), .Cin(s1_310_hacout), .S(s2_327_fas), .Cout(s2_327_facout));
full_adder s2_32fa8 ( .A(s1_320_fas), .B(s1_321_fas), .Cin(s1_322_fas), .S(s2_328_fas), .Cout(s2_328_facout));
full_adder s2_33fa0 ( .A(ps_3322), .B(ps_3321), .Cin(ps_3320), .S(s2_330_fas), .Cout(s2_330_facout));
full_adder s2_33fa1 ( .A(ps_3319), .B(ps_3318), .Cin(ps_3317), .S(s2_331_fas), .Cout(s2_331_facout));
full_adder s2_33fa2 ( .A(ps_3316), .B(ps_3315), .Cin(ps_3314), .S(s2_332_fas), .Cout(s2_332_facout));
full_adder s2_33fa3 ( .A(ps_3313), .B(ps_3312), .Cin(ps_3311), .S(s2_333_fas), .Cout(s2_333_facout));
full_adder s2_33fa4 ( .A(ps_3310), .B(ps_339), .Cin(ps_338), .S(s2_334_fas), .Cout(s2_334_facout));
full_adder s2_33fa5 ( .A(ps_337), .B(ps_336), .Cin(ps_335), .S(s2_335_fas), .Cout(s2_335_facout));
full_adder s2_33fa6 ( .A(ps_334), .B(ps_333), .Cin(ps_332), .S(s2_336_fas), .Cout(s2_336_facout));
full_adder s2_33fa7 ( .A(s1_320_facout), .B(s1_321_facout), .Cin(s1_322_facout), .S(s2_337_fas), .Cout(s2_337_facout));
full_adder s2_33fa8 ( .A(s1_320_hacout), .B(s1_330_fas), .Cin(s1_331_fas), .S(s2_338_fas), .Cout(s2_338_facout));
full_adder s2_34fa0 ( .A(ps_3425), .B(ps_3424), .Cin(ps_3423), .S(s2_340_fas), .Cout(s2_340_facout));
full_adder s2_34fa1 ( .A(ps_3422), .B(ps_3421), .Cin(ps_3420), .S(s2_341_fas), .Cout(s2_341_facout));
full_adder s2_34fa2 ( .A(ps_3419), .B(ps_3418), .Cin(ps_3417), .S(s2_342_fas), .Cout(s2_342_facout));
full_adder s2_34fa3 ( .A(ps_3416), .B(ps_3415), .Cin(ps_3414), .S(s2_343_fas), .Cout(s2_343_facout));
full_adder s2_34fa4 ( .A(ps_3413), .B(ps_3412), .Cin(ps_3411), .S(s2_344_fas), .Cout(s2_344_facout));
full_adder s2_34fa5 ( .A(ps_3410), .B(ps_349), .Cin(ps_348), .S(s2_345_fas), .Cout(s2_345_facout));
full_adder s2_34fa6 ( .A(ps_347), .B(ps_346), .Cin(ps_345), .S(s2_346_fas), .Cout(s2_346_facout));
full_adder s2_34fa7 ( .A(ps_344), .B(ps_343), .Cin(s1_330_facout), .S(s2_347_fas), .Cout(s2_347_facout));
full_adder s2_34fa8 ( .A(s1_331_facout), .B(s1_332_facout), .Cin(s1_340_fas), .S(s2_348_fas), .Cout(s2_348_facout));
full_adder s2_35fa0 ( .A(ps_3528), .B(ps_3527), .Cin(ps_3526), .S(s2_350_fas), .Cout(s2_350_facout));
full_adder s2_35fa1 ( .A(ps_3525), .B(ps_3524), .Cin(ps_3523), .S(s2_351_fas), .Cout(s2_351_facout));
full_adder s2_35fa2 ( .A(ps_3522), .B(ps_3521), .Cin(ps_3520), .S(s2_352_fas), .Cout(s2_352_facout));
full_adder s2_35fa3 ( .A(ps_3519), .B(ps_3518), .Cin(ps_3517), .S(s2_353_fas), .Cout(s2_353_facout));
full_adder s2_35fa4 ( .A(ps_3516), .B(ps_3515), .Cin(ps_3514), .S(s2_354_fas), .Cout(s2_354_facout));
full_adder s2_35fa5 ( .A(ps_3513), .B(ps_3512), .Cin(ps_3511), .S(s2_355_fas), .Cout(s2_355_facout));
full_adder s2_35fa6 ( .A(ps_3510), .B(ps_359), .Cin(ps_358), .S(s2_356_fas), .Cout(s2_356_facout));
full_adder s2_35fa7 ( .A(ps_357), .B(ps_356), .Cin(ps_355), .S(s2_357_fas), .Cout(s2_357_facout));
full_adder s2_35fa8 ( .A(ps_354), .B(s1_340_facout), .Cin(s1_341_facout), .S(s2_358_fas), .Cout(s2_358_facout));
full_adder s2_36fa0 ( .A(ps_3631), .B(ps_3630), .Cin(ps_3629), .S(s2_360_fas), .Cout(s2_360_facout));
full_adder s2_36fa1 ( .A(ps_3628), .B(ps_3627), .Cin(ps_3626), .S(s2_361_fas), .Cout(s2_361_facout));
full_adder s2_36fa2 ( .A(ps_3625), .B(ps_3624), .Cin(ps_3623), .S(s2_362_fas), .Cout(s2_362_facout));
full_adder s2_36fa3 ( .A(ps_3622), .B(ps_3621), .Cin(ps_3620), .S(s2_363_fas), .Cout(s2_363_facout));
full_adder s2_36fa4 ( .A(ps_3619), .B(ps_3618), .Cin(ps_3617), .S(s2_364_fas), .Cout(s2_364_facout));
full_adder s2_36fa5 ( .A(ps_3616), .B(ps_3615), .Cin(ps_3614), .S(s2_365_fas), .Cout(s2_365_facout));
full_adder s2_36fa6 ( .A(ps_3613), .B(ps_3612), .Cin(ps_3611), .S(s2_366_fas), .Cout(s2_366_facout));
full_adder s2_36fa7 ( .A(ps_3610), .B(ps_369), .Cin(ps_368), .S(s2_367_fas), .Cout(s2_367_facout));
full_adder s2_36fa8 ( .A(ps_367), .B(ps_366), .Cin(ps_365), .S(s2_368_fas), .Cout(s2_368_facout));
full_adder s2_37fa0 ( .A(ps_3731), .B(ps_3730), .Cin(ps_3729), .S(s2_370_fas), .Cout(s2_370_facout));
full_adder s2_37fa1 ( .A(ps_3728), .B(ps_3727), .Cin(ps_3726), .S(s2_371_fas), .Cout(s2_371_facout));
full_adder s2_37fa2 ( .A(ps_3725), .B(ps_3724), .Cin(ps_3723), .S(s2_372_fas), .Cout(s2_372_facout));
full_adder s2_37fa3 ( .A(ps_3722), .B(ps_3721), .Cin(ps_3720), .S(s2_373_fas), .Cout(s2_373_facout));
full_adder s2_37fa4 ( .A(ps_3719), .B(ps_3718), .Cin(ps_3717), .S(s2_374_fas), .Cout(s2_374_facout));
full_adder s2_37fa5 ( .A(ps_3716), .B(ps_3715), .Cin(ps_3714), .S(s2_375_fas), .Cout(s2_375_facout));
full_adder s2_37fa6 ( .A(ps_3713), .B(ps_3712), .Cin(ps_3711), .S(s2_376_fas), .Cout(s2_376_facout));
full_adder s2_37fa7 ( .A(ps_3710), .B(ps_379), .Cin(ps_378), .S(s2_377_fas), .Cout(s2_377_facout));
full_adder s2_38fa0 ( .A(ps_3831), .B(ps_3830), .Cin(ps_3829), .S(s2_380_fas), .Cout(s2_380_facout));
full_adder s2_38fa1 ( .A(ps_3828), .B(ps_3827), .Cin(ps_3826), .S(s2_381_fas), .Cout(s2_381_facout));
full_adder s2_38fa2 ( .A(ps_3825), .B(ps_3824), .Cin(ps_3823), .S(s2_382_fas), .Cout(s2_382_facout));
full_adder s2_38fa3 ( .A(ps_3822), .B(ps_3821), .Cin(ps_3820), .S(s2_383_fas), .Cout(s2_383_facout));
full_adder s2_38fa4 ( .A(ps_3819), .B(ps_3818), .Cin(ps_3817), .S(s2_384_fas), .Cout(s2_384_facout));
full_adder s2_38fa5 ( .A(ps_3816), .B(ps_3815), .Cin(ps_3814), .S(s2_385_fas), .Cout(s2_385_facout));
full_adder s2_38fa6 ( .A(ps_3813), .B(ps_3812), .Cin(ps_3811), .S(s2_386_fas), .Cout(s2_386_facout));
full_adder s2_39fa0 ( .A(ps_3931), .B(ps_3930), .Cin(ps_3929), .S(s2_390_fas), .Cout(s2_390_facout));
full_adder s2_39fa1 ( .A(ps_3928), .B(ps_3927), .Cin(ps_3926), .S(s2_391_fas), .Cout(s2_391_facout));
full_adder s2_39fa2 ( .A(ps_3925), .B(ps_3924), .Cin(ps_3923), .S(s2_392_fas), .Cout(s2_392_facout));
full_adder s2_39fa3 ( .A(ps_3922), .B(ps_3921), .Cin(ps_3920), .S(s2_393_fas), .Cout(s2_393_facout));
full_adder s2_39fa4 ( .A(ps_3919), .B(ps_3918), .Cin(ps_3917), .S(s2_394_fas), .Cout(s2_394_facout));
full_adder s2_39fa5 ( .A(ps_3916), .B(ps_3915), .Cin(ps_3914), .S(s2_395_fas), .Cout(s2_395_facout));
full_adder s2_40fa0 ( .A(ps_4031), .B(ps_4030), .Cin(ps_4029), .S(s2_400_fas), .Cout(s2_400_facout));
full_adder s2_40fa1 ( .A(ps_4028), .B(ps_4027), .Cin(ps_4026), .S(s2_401_fas), .Cout(s2_401_facout));
full_adder s2_40fa2 ( .A(ps_4025), .B(ps_4024), .Cin(ps_4023), .S(s2_402_fas), .Cout(s2_402_facout));
full_adder s2_40fa3 ( .A(ps_4022), .B(ps_4021), .Cin(ps_4020), .S(s2_403_fas), .Cout(s2_403_facout));
full_adder s2_40fa4 ( .A(ps_4019), .B(ps_4018), .Cin(ps_4017), .S(s2_404_fas), .Cout(s2_404_facout));
full_adder s2_41fa0 ( .A(ps_4131), .B(ps_4130), .Cin(ps_4129), .S(s2_410_fas), .Cout(s2_410_facout));
full_adder s2_41fa1 ( .A(ps_4128), .B(ps_4127), .Cin(ps_4126), .S(s2_411_fas), .Cout(s2_411_facout));
full_adder s2_41fa2 ( .A(ps_4125), .B(ps_4124), .Cin(ps_4123), .S(s2_412_fas), .Cout(s2_412_facout));
full_adder s2_41fa3 ( .A(ps_4122), .B(ps_4121), .Cin(ps_4120), .S(s2_413_fas), .Cout(s2_413_facout));
full_adder s2_42fa0 ( .A(ps_4231), .B(ps_4230), .Cin(ps_4229), .S(s2_420_fas), .Cout(s2_420_facout));
full_adder s2_42fa1 ( .A(ps_4228), .B(ps_4227), .Cin(ps_4226), .S(s2_421_fas), .Cout(s2_421_facout));
full_adder s2_42fa2 ( .A(ps_4225), .B(ps_4224), .Cin(ps_4223), .S(s2_422_fas), .Cout(s2_422_facout));
full_adder s2_43fa0 ( .A(ps_4331), .B(ps_4330), .Cin(ps_4329), .S(s2_430_fas), .Cout(s2_430_facout));
full_adder s2_43fa1 ( .A(ps_4328), .B(ps_4327), .Cin(ps_4326), .S(s2_431_fas), .Cout(s2_431_facout));
full_adder s2_44fa0 ( .A(ps_4431), .B(ps_4430), .Cin(ps_4429), .S(s2_440_fas), .Cout(s2_440_facout));
logic s3_130_hacout, s3_130_has, s3_140_facout, s3_140_fas, s3_140_hacout, s3_140_has, s3_150_facout, s3_150_fas, s3_151_facout, s3_151_fas, s3_150_hacout, s3_150_has, s3_160_facout, s3_160_fas, s3_161_facout, s3_161_fas, s3_162_facout, s3_162_fas, s3_160_hacout, s3_160_has, s3_170_facout, s3_170_fas, s3_171_facout, s3_171_fas, s3_172_facout, s3_172_fas, s3_173_facout, s3_173_fas, s3_170_hacout, s3_170_has, s3_180_facout, s3_180_fas, s3_181_facout, s3_181_fas, s3_182_facout, s3_182_fas, s3_183_facout, s3_183_fas, s3_184_facout, s3_184_fas, s3_180_hacout, s3_180_has, s3_190_facout, s3_190_fas, s3_191_facout, s3_191_fas, s3_192_facout, s3_192_fas, s3_193_facout, s3_193_fas, s3_194_facout, s3_194_fas, s3_195_facout, s3_195_fas, s3_200_facout, s3_200_fas, s3_201_facout, s3_201_fas, s3_202_facout, s3_202_fas, s3_203_facout, s3_203_fas, s3_204_facout, s3_204_fas, s3_205_facout, s3_205_fas, s3_210_facout, s3_210_fas, s3_211_facout, s3_211_fas, s3_212_facout, s3_212_fas, s3_213_facout, s3_213_fas, s3_214_facout, s3_214_fas, s3_215_facout, s3_215_fas, s3_220_facout, s3_220_fas, s3_221_facout, s3_221_fas, s3_222_facout, s3_222_fas, s3_223_facout, s3_223_fas, s3_224_facout, s3_224_fas, s3_225_facout, s3_225_fas, s3_230_facout, s3_230_fas, s3_231_facout, s3_231_fas, s3_232_facout, s3_232_fas, s3_233_facout, s3_233_fas, s3_234_facout, s3_234_fas, s3_235_facout, s3_235_fas, s3_240_facout, s3_240_fas, s3_241_facout, s3_241_fas, s3_242_facout, s3_242_fas, s3_243_facout, s3_243_fas, s3_244_facout, s3_244_fas, s3_245_facout, s3_245_fas, s3_250_facout, s3_250_fas, s3_251_facout, s3_251_fas, s3_252_facout, s3_252_fas, s3_253_facout, s3_253_fas, s3_254_facout, s3_254_fas, s3_255_facout, s3_255_fas, s3_260_facout, s3_260_fas, s3_261_facout, s3_261_fas, s3_262_facout, s3_262_fas, s3_263_facout, s3_263_fas, s3_264_facout, s3_264_fas, s3_265_facout, s3_265_fas, s3_270_facout, s3_270_fas, s3_271_facout, s3_271_fas, s3_272_facout, s3_272_fas, s3_273_facout, s3_273_fas, s3_274_facout, s3_274_fas, s3_275_facout, s3_275_fas, s3_280_facout, s3_280_fas, s3_281_facout, s3_281_fas, s3_282_facout, s3_282_fas, s3_283_facout, s3_283_fas, s3_284_facout, s3_284_fas, s3_285_facout, s3_285_fas, s3_290_facout, s3_290_fas, s3_291_facout, s3_291_fas, s3_292_facout, s3_292_fas, s3_293_facout, s3_293_fas, s3_294_facout, s3_294_fas, s3_295_facout, s3_295_fas, s3_300_facout, s3_300_fas, s3_301_facout, s3_301_fas, s3_302_facout, s3_302_fas, s3_303_facout, s3_303_fas, s3_304_facout, s3_304_fas, s3_305_facout, s3_305_fas, s3_310_facout, s3_310_fas, s3_311_facout, s3_311_fas, s3_312_facout, s3_312_fas, s3_313_facout, s3_313_fas, s3_314_facout, s3_314_fas, s3_315_facout, s3_315_fas, s3_320_facout, s3_320_fas, s3_321_facout, s3_321_fas, s3_322_facout, s3_322_fas, s3_323_facout, s3_323_fas, s3_324_facout, s3_324_fas, s3_325_facout, s3_325_fas, s3_330_facout, s3_330_fas, s3_331_facout, s3_331_fas, s3_332_facout, s3_332_fas, s3_333_facout, s3_333_fas, s3_334_facout, s3_334_fas, s3_335_facout, s3_335_fas, s3_340_facout, s3_340_fas, s3_341_facout, s3_341_fas, s3_342_facout, s3_342_fas, s3_343_facout, s3_343_fas, s3_344_facout, s3_344_fas, s3_345_facout, s3_345_fas, s3_350_facout, s3_350_fas, s3_351_facout, s3_351_fas, s3_352_facout, s3_352_fas, s3_353_facout, s3_353_fas, s3_354_facout, s3_354_fas, s3_355_facout, s3_355_fas, s3_360_facout, s3_360_fas, s3_361_facout, s3_361_fas, s3_362_facout, s3_362_fas, s3_363_facout, s3_363_fas, s3_364_facout, s3_364_fas, s3_365_facout, s3_365_fas, s3_370_facout, s3_370_fas, s3_371_facout, s3_371_fas, s3_372_facout, s3_372_fas, s3_373_facout, s3_373_fas, s3_374_facout, s3_374_fas, s3_375_facout, s3_375_fas, s3_380_facout, s3_380_fas, s3_381_facout, s3_381_fas, s3_382_facout, s3_382_fas, s3_383_facout, s3_383_fas, s3_384_facout, s3_384_fas, s3_385_facout, s3_385_fas, s3_390_facout, s3_390_fas, s3_391_facout, s3_391_fas, s3_392_facout, s3_392_fas, s3_393_facout, s3_393_fas, s3_394_facout, s3_394_fas, s3_395_facout, s3_395_fas, s3_400_facout, s3_400_fas, s3_401_facout, s3_401_fas, s3_402_facout, s3_402_fas, s3_403_facout, s3_403_fas, s3_404_facout, s3_404_fas, s3_405_facout, s3_405_fas, s3_410_facout, s3_410_fas, s3_411_facout, s3_411_fas, s3_412_facout, s3_412_fas, s3_413_facout, s3_413_fas, s3_414_facout, s3_414_fas, s3_415_facout, s3_415_fas, s3_420_facout, s3_420_fas, s3_421_facout, s3_421_fas, s3_422_facout, s3_422_fas, s3_423_facout, s3_423_fas, s3_424_facout, s3_424_fas, s3_425_facout, s3_425_fas, s3_430_facout, s3_430_fas, s3_431_facout, s3_431_fas, s3_432_facout, s3_432_fas, s3_433_facout, s3_433_fas, s3_434_facout, s3_434_fas, s3_435_facout, s3_435_fas, s3_440_facout, s3_440_fas, s3_441_facout, s3_441_fas, s3_442_facout, s3_442_fas, s3_443_facout, s3_443_fas, s3_444_facout, s3_444_fas, s3_445_facout, s3_445_fas, s3_450_facout, s3_450_fas, s3_451_facout, s3_451_fas, s3_452_facout, s3_452_fas, s3_453_facout, s3_453_fas, s3_454_facout, s3_454_fas, s3_455_facout, s3_455_fas, s3_460_facout, s3_460_fas, s3_461_facout, s3_461_fas, s3_462_facout, s3_462_fas, s3_463_facout, s3_463_fas, s3_464_facout, s3_464_fas, s3_470_facout, s3_470_fas, s3_471_facout, s3_471_fas, s3_472_facout, s3_472_fas, s3_473_facout, s3_473_fas, s3_480_facout, s3_480_fas, s3_481_facout, s3_481_fas, s3_482_facout, s3_482_fas, s3_490_facout, s3_490_fas, s3_491_facout, s3_491_fas, s3_500_facout, s3_500_fas;
/* ========================= Stage 3 ========================= */
half_adder s3_13ha0 ( .A(ps_1313), .B(ps_1312), .S(s3_130_has), .Cout(s3_130_hacout));
full_adder s3_14fa0 ( .A(ps_1414), .B(ps_1413), .Cin(ps_1412), .S(s3_140_fas), .Cout(s3_140_facout));
half_adder s3_14ha0 ( .A(ps_1411), .B(ps_1410), .S(s3_140_has), .Cout(s3_140_hacout));
full_adder s3_15fa0 ( .A(ps_1515), .B(ps_1514), .Cin(ps_1513), .S(s3_150_fas), .Cout(s3_150_facout));
full_adder s3_15fa1 ( .A(ps_1512), .B(ps_1511), .Cin(ps_1510), .S(s3_151_fas), .Cout(s3_151_facout));
half_adder s3_15ha0 ( .A(ps_159), .B(ps_158), .S(s3_150_has), .Cout(s3_150_hacout));
full_adder s3_16fa0 ( .A(ps_1616), .B(ps_1615), .Cin(ps_1614), .S(s3_160_fas), .Cout(s3_160_facout));
full_adder s3_16fa1 ( .A(ps_1613), .B(ps_1612), .Cin(ps_1611), .S(s3_161_fas), .Cout(s3_161_facout));
full_adder s3_16fa2 ( .A(ps_1610), .B(ps_169), .Cin(ps_168), .S(s3_162_fas), .Cout(s3_162_facout));
half_adder s3_16ha0 ( .A(ps_167), .B(ps_166), .S(s3_160_has), .Cout(s3_160_hacout));
full_adder s3_17fa0 ( .A(ps_1717), .B(ps_1716), .Cin(ps_1715), .S(s3_170_fas), .Cout(s3_170_facout));
full_adder s3_17fa1 ( .A(ps_1714), .B(ps_1713), .Cin(ps_1712), .S(s3_171_fas), .Cout(s3_171_facout));
full_adder s3_17fa2 ( .A(ps_1711), .B(ps_1710), .Cin(ps_179), .S(s3_172_fas), .Cout(s3_172_facout));
full_adder s3_17fa3 ( .A(ps_178), .B(ps_177), .Cin(ps_176), .S(s3_173_fas), .Cout(s3_173_facout));
half_adder s3_17ha0 ( .A(ps_175), .B(ps_174), .S(s3_170_has), .Cout(s3_170_hacout));
full_adder s3_18fa0 ( .A(ps_1818), .B(ps_1817), .Cin(ps_1816), .S(s3_180_fas), .Cout(s3_180_facout));
full_adder s3_18fa1 ( .A(ps_1815), .B(ps_1814), .Cin(ps_1813), .S(s3_181_fas), .Cout(s3_181_facout));
full_adder s3_18fa2 ( .A(ps_1812), .B(ps_1811), .Cin(ps_1810), .S(s3_182_fas), .Cout(s3_182_facout));
full_adder s3_18fa3 ( .A(ps_189), .B(ps_188), .Cin(ps_187), .S(s3_183_fas), .Cout(s3_183_facout));
full_adder s3_18fa4 ( .A(ps_186), .B(ps_185), .Cin(ps_184), .S(s3_184_fas), .Cout(s3_184_facout));
half_adder s3_18ha0 ( .A(ps_183), .B(ps_182), .S(s3_180_has), .Cout(s3_180_hacout));
full_adder s3_19fa0 ( .A(ps_1917), .B(ps_1916), .Cin(ps_1915), .S(s3_190_fas), .Cout(s3_190_facout));
full_adder s3_19fa1 ( .A(ps_1914), .B(ps_1913), .Cin(ps_1912), .S(s3_191_fas), .Cout(s3_191_facout));
full_adder s3_19fa2 ( .A(ps_1911), .B(ps_1910), .Cin(ps_199), .S(s3_192_fas), .Cout(s3_192_facout));
full_adder s3_19fa3 ( .A(ps_198), .B(ps_197), .Cin(ps_196), .S(s3_193_fas), .Cout(s3_193_facout));
full_adder s3_19fa4 ( .A(ps_195), .B(ps_194), .Cin(ps_193), .S(s3_194_fas), .Cout(s3_194_facout));
full_adder s3_19fa5 ( .A(ps_192), .B(ps_191), .Cin(ps_190), .S(s3_195_fas), .Cout(s3_195_facout));
full_adder s3_20fa0 ( .A(ps_2015), .B(ps_2014), .Cin(ps_2013), .S(s3_200_fas), .Cout(s3_200_facout));
full_adder s3_20fa1 ( .A(ps_2012), .B(ps_2011), .Cin(ps_2010), .S(s3_201_fas), .Cout(s3_201_facout));
full_adder s3_20fa2 ( .A(ps_209), .B(ps_208), .Cin(ps_207), .S(s3_202_fas), .Cout(s3_202_facout));
full_adder s3_20fa3 ( .A(ps_206), .B(ps_205), .Cin(ps_204), .S(s3_203_fas), .Cout(s3_203_facout));
full_adder s3_20fa4 ( .A(ps_203), .B(ps_202), .Cin(ps_201), .S(s3_204_fas), .Cout(s3_204_facout));
full_adder s3_20fa5 ( .A(ps_200), .B(s2_190_hacout), .Cin(s2_200_fas), .S(s3_205_fas), .Cout(s3_205_facout));
full_adder s3_21fa0 ( .A(ps_2113), .B(ps_2112), .Cin(ps_2111), .S(s3_210_fas), .Cout(s3_210_facout));
full_adder s3_21fa1 ( .A(ps_2110), .B(ps_219), .Cin(ps_218), .S(s3_211_fas), .Cout(s3_211_facout));
full_adder s3_21fa2 ( .A(ps_217), .B(ps_216), .Cin(ps_215), .S(s3_212_fas), .Cout(s3_212_facout));
full_adder s3_21fa3 ( .A(ps_214), .B(ps_213), .Cin(ps_212), .S(s3_213_fas), .Cout(s3_213_facout));
full_adder s3_21fa4 ( .A(ps_211), .B(ps_210), .Cin(s2_200_facout), .S(s3_214_fas), .Cout(s3_214_facout));
full_adder s3_21fa5 ( .A(s2_200_hacout), .B(s2_210_fas), .Cin(s2_211_fas), .S(s3_215_fas), .Cout(s3_215_facout));
full_adder s3_22fa0 ( .A(ps_2211), .B(ps_2210), .Cin(ps_229), .S(s3_220_fas), .Cout(s3_220_facout));
full_adder s3_22fa1 ( .A(ps_228), .B(ps_227), .Cin(ps_226), .S(s3_221_fas), .Cout(s3_221_facout));
full_adder s3_22fa2 ( .A(ps_225), .B(ps_224), .Cin(ps_223), .S(s3_222_fas), .Cout(s3_222_facout));
full_adder s3_22fa3 ( .A(ps_222), .B(ps_221), .Cin(ps_220), .S(s3_223_fas), .Cout(s3_223_facout));
full_adder s3_22fa4 ( .A(s2_210_facout), .B(s2_211_facout), .Cin(s2_210_hacout), .S(s3_224_fas), .Cout(s3_224_facout));
full_adder s3_22fa5 ( .A(s2_220_fas), .B(s2_221_fas), .Cin(s2_222_fas), .S(s3_225_fas), .Cout(s3_225_facout));
full_adder s3_23fa0 ( .A(ps_239), .B(ps_238), .Cin(ps_237), .S(s3_230_fas), .Cout(s3_230_facout));
full_adder s3_23fa1 ( .A(ps_236), .B(ps_235), .Cin(ps_234), .S(s3_231_fas), .Cout(s3_231_facout));
full_adder s3_23fa2 ( .A(ps_233), .B(ps_232), .Cin(ps_231), .S(s3_232_fas), .Cout(s3_232_facout));
full_adder s3_23fa3 ( .A(ps_230), .B(s2_220_facout), .Cin(s2_221_facout), .S(s3_233_fas), .Cout(s3_233_facout));
full_adder s3_23fa4 ( .A(s2_222_facout), .B(s2_220_hacout), .Cin(s2_230_fas), .S(s3_234_fas), .Cout(s3_234_facout));
full_adder s3_23fa5 ( .A(s2_231_fas), .B(s2_232_fas), .Cin(s2_233_fas), .S(s3_235_fas), .Cout(s3_235_facout));
full_adder s3_24fa0 ( .A(ps_247), .B(ps_246), .Cin(ps_245), .S(s3_240_fas), .Cout(s3_240_facout));
full_adder s3_24fa1 ( .A(ps_244), .B(ps_243), .Cin(ps_242), .S(s3_241_fas), .Cout(s3_241_facout));
full_adder s3_24fa2 ( .A(ps_241), .B(ps_240), .Cin(s2_230_facout), .S(s3_242_fas), .Cout(s3_242_facout));
full_adder s3_24fa3 ( .A(s2_231_facout), .B(s2_232_facout), .Cin(s2_233_facout), .S(s3_243_fas), .Cout(s3_243_facout));
full_adder s3_24fa4 ( .A(s2_230_hacout), .B(s2_240_fas), .Cin(s2_241_fas), .S(s3_244_fas), .Cout(s3_244_facout));
full_adder s3_24fa5 ( .A(s2_242_fas), .B(s2_243_fas), .Cin(s2_244_fas), .S(s3_245_fas), .Cout(s3_245_facout));
full_adder s3_25fa0 ( .A(ps_255), .B(ps_254), .Cin(ps_253), .S(s3_250_fas), .Cout(s3_250_facout));
full_adder s3_25fa1 ( .A(ps_252), .B(ps_251), .Cin(ps_250), .S(s3_251_fas), .Cout(s3_251_facout));
full_adder s3_25fa2 ( .A(s2_240_facout), .B(s2_241_facout), .Cin(s2_242_facout), .S(s3_252_fas), .Cout(s3_252_facout));
full_adder s3_25fa3 ( .A(s2_243_facout), .B(s2_244_facout), .Cin(s2_240_hacout), .S(s3_253_fas), .Cout(s3_253_facout));
full_adder s3_25fa4 ( .A(s2_250_fas), .B(s2_251_fas), .Cin(s2_252_fas), .S(s3_254_fas), .Cout(s3_254_facout));
full_adder s3_25fa5 ( .A(s2_253_fas), .B(s2_254_fas), .Cin(s2_255_fas), .S(s3_255_fas), .Cout(s3_255_facout));
full_adder s3_26fa0 ( .A(ps_263), .B(ps_262), .Cin(ps_261), .S(s3_260_fas), .Cout(s3_260_facout));
full_adder s3_26fa1 ( .A(ps_260), .B(s2_250_facout), .Cin(s2_251_facout), .S(s3_261_fas), .Cout(s3_261_facout));
full_adder s3_26fa2 ( .A(s2_252_facout), .B(s2_253_facout), .Cin(s2_254_facout), .S(s3_262_fas), .Cout(s3_262_facout));
full_adder s3_26fa3 ( .A(s2_255_facout), .B(s2_250_hacout), .Cin(s2_260_fas), .S(s3_263_fas), .Cout(s3_263_facout));
full_adder s3_26fa4 ( .A(s2_261_fas), .B(s2_262_fas), .Cin(s2_263_fas), .S(s3_264_fas), .Cout(s3_264_facout));
full_adder s3_26fa5 ( .A(s2_264_fas), .B(s2_265_fas), .Cin(s2_266_fas), .S(s3_265_fas), .Cout(s3_265_facout));
full_adder s3_27fa0 ( .A(ps_271), .B(ps_270), .Cin(s2_260_facout), .S(s3_270_fas), .Cout(s3_270_facout));
full_adder s3_27fa1 ( .A(s2_261_facout), .B(s2_262_facout), .Cin(s2_263_facout), .S(s3_271_fas), .Cout(s3_271_facout));
full_adder s3_27fa2 ( .A(s2_264_facout), .B(s2_265_facout), .Cin(s2_266_facout), .S(s3_272_fas), .Cout(s3_272_facout));
full_adder s3_27fa3 ( .A(s2_260_hacout), .B(s2_270_fas), .Cin(s2_271_fas), .S(s3_273_fas), .Cout(s3_273_facout));
full_adder s3_27fa4 ( .A(s2_272_fas), .B(s2_273_fas), .Cin(s2_274_fas), .S(s3_274_fas), .Cout(s3_274_facout));
full_adder s3_27fa5 ( .A(s2_275_fas), .B(s2_276_fas), .Cin(s2_277_fas), .S(s3_275_fas), .Cout(s3_275_facout));
full_adder s3_28fa0 ( .A(s1_280_has), .B(s2_270_facout), .Cin(s2_271_facout), .S(s3_280_fas), .Cout(s3_280_facout));
full_adder s3_28fa1 ( .A(s2_272_facout), .B(s2_273_facout), .Cin(s2_274_facout), .S(s3_281_fas), .Cout(s3_281_facout));
full_adder s3_28fa2 ( .A(s2_275_facout), .B(s2_276_facout), .Cin(s2_277_facout), .S(s3_282_fas), .Cout(s3_282_facout));
full_adder s3_28fa3 ( .A(s2_270_hacout), .B(s2_280_fas), .Cin(s2_281_fas), .S(s3_283_fas), .Cout(s3_283_facout));
full_adder s3_28fa4 ( .A(s2_282_fas), .B(s2_283_fas), .Cin(s2_284_fas), .S(s3_284_fas), .Cout(s3_284_facout));
full_adder s3_28fa5 ( .A(s2_285_fas), .B(s2_286_fas), .Cin(s2_287_fas), .S(s3_285_fas), .Cout(s3_285_facout));
full_adder s3_29fa0 ( .A(s1_290_has), .B(s2_280_facout), .Cin(s2_281_facout), .S(s3_290_fas), .Cout(s3_290_facout));
full_adder s3_29fa1 ( .A(s2_282_facout), .B(s2_283_facout), .Cin(s2_284_facout), .S(s3_291_fas), .Cout(s3_291_facout));
full_adder s3_29fa2 ( .A(s2_285_facout), .B(s2_286_facout), .Cin(s2_287_facout), .S(s3_292_fas), .Cout(s3_292_facout));
full_adder s3_29fa3 ( .A(s2_288_facout), .B(s2_290_fas), .Cin(s2_291_fas), .S(s3_293_fas), .Cout(s3_293_facout));
full_adder s3_29fa4 ( .A(s2_292_fas), .B(s2_293_fas), .Cin(s2_294_fas), .S(s3_294_fas), .Cout(s3_294_facout));
full_adder s3_29fa5 ( .A(s2_295_fas), .B(s2_296_fas), .Cin(s2_297_fas), .S(s3_295_fas), .Cout(s3_295_facout));
full_adder s3_30fa0 ( .A(s1_300_has), .B(s2_290_facout), .Cin(s2_291_facout), .S(s3_300_fas), .Cout(s3_300_facout));
full_adder s3_30fa1 ( .A(s2_292_facout), .B(s2_293_facout), .Cin(s2_294_facout), .S(s3_301_fas), .Cout(s3_301_facout));
full_adder s3_30fa2 ( .A(s2_295_facout), .B(s2_296_facout), .Cin(s2_297_facout), .S(s3_302_fas), .Cout(s3_302_facout));
full_adder s3_30fa3 ( .A(s2_298_facout), .B(s2_300_fas), .Cin(s2_301_fas), .S(s3_303_fas), .Cout(s3_303_facout));
full_adder s3_30fa4 ( .A(s2_302_fas), .B(s2_303_fas), .Cin(s2_304_fas), .S(s3_304_fas), .Cout(s3_304_facout));
full_adder s3_30fa5 ( .A(s2_305_fas), .B(s2_306_fas), .Cin(s2_307_fas), .S(s3_305_fas), .Cout(s3_305_facout));
full_adder s3_31fa0 ( .A(s1_310_has), .B(s2_300_facout), .Cin(s2_301_facout), .S(s3_310_fas), .Cout(s3_310_facout));
full_adder s3_31fa1 ( .A(s2_302_facout), .B(s2_303_facout), .Cin(s2_304_facout), .S(s3_311_fas), .Cout(s3_311_facout));
full_adder s3_31fa2 ( .A(s2_305_facout), .B(s2_306_facout), .Cin(s2_307_facout), .S(s3_312_fas), .Cout(s3_312_facout));
full_adder s3_31fa3 ( .A(s2_308_facout), .B(s2_310_fas), .Cin(s2_311_fas), .S(s3_313_fas), .Cout(s3_313_facout));
full_adder s3_31fa4 ( .A(s2_312_fas), .B(s2_313_fas), .Cin(s2_314_fas), .S(s3_314_fas), .Cout(s3_314_facout));
full_adder s3_31fa5 ( .A(s2_315_fas), .B(s2_316_fas), .Cin(s2_317_fas), .S(s3_315_fas), .Cout(s3_315_facout));
full_adder s3_32fa0 ( .A(s1_320_has), .B(s2_310_facout), .Cin(s2_311_facout), .S(s3_320_fas), .Cout(s3_320_facout));
full_adder s3_32fa1 ( .A(s2_312_facout), .B(s2_313_facout), .Cin(s2_314_facout), .S(s3_321_fas), .Cout(s3_321_facout));
full_adder s3_32fa2 ( .A(s2_315_facout), .B(s2_316_facout), .Cin(s2_317_facout), .S(s3_322_fas), .Cout(s3_322_facout));
full_adder s3_32fa3 ( .A(s2_318_facout), .B(s2_320_fas), .Cin(s2_321_fas), .S(s3_323_fas), .Cout(s3_323_facout));
full_adder s3_32fa4 ( .A(s2_322_fas), .B(s2_323_fas), .Cin(s2_324_fas), .S(s3_324_fas), .Cout(s3_324_facout));
full_adder s3_32fa5 ( .A(s2_325_fas), .B(s2_326_fas), .Cin(s2_327_fas), .S(s3_325_fas), .Cout(s3_325_facout));
full_adder s3_33fa0 ( .A(s1_332_fas), .B(s2_320_facout), .Cin(s2_321_facout), .S(s3_330_fas), .Cout(s3_330_facout));
full_adder s3_33fa1 ( .A(s2_322_facout), .B(s2_323_facout), .Cin(s2_324_facout), .S(s3_331_fas), .Cout(s3_331_facout));
full_adder s3_33fa2 ( .A(s2_325_facout), .B(s2_326_facout), .Cin(s2_327_facout), .S(s3_332_fas), .Cout(s3_332_facout));
full_adder s3_33fa3 ( .A(s2_328_facout), .B(s2_330_fas), .Cin(s2_331_fas), .S(s3_333_fas), .Cout(s3_333_facout));
full_adder s3_33fa4 ( .A(s2_332_fas), .B(s2_333_fas), .Cin(s2_334_fas), .S(s3_334_fas), .Cout(s3_334_facout));
full_adder s3_33fa5 ( .A(s2_335_fas), .B(s2_336_fas), .Cin(s2_337_fas), .S(s3_335_fas), .Cout(s3_335_facout));
full_adder s3_34fa0 ( .A(s1_341_fas), .B(s2_330_facout), .Cin(s2_331_facout), .S(s3_340_fas), .Cout(s3_340_facout));
full_adder s3_34fa1 ( .A(s2_332_facout), .B(s2_333_facout), .Cin(s2_334_facout), .S(s3_341_fas), .Cout(s3_341_facout));
full_adder s3_34fa2 ( .A(s2_335_facout), .B(s2_336_facout), .Cin(s2_337_facout), .S(s3_342_fas), .Cout(s3_342_facout));
full_adder s3_34fa3 ( .A(s2_338_facout), .B(s2_340_fas), .Cin(s2_341_fas), .S(s3_343_fas), .Cout(s3_343_facout));
full_adder s3_34fa4 ( .A(s2_342_fas), .B(s2_343_fas), .Cin(s2_344_fas), .S(s3_344_fas), .Cout(s3_344_facout));
full_adder s3_34fa5 ( .A(s2_345_fas), .B(s2_346_fas), .Cin(s2_347_fas), .S(s3_345_fas), .Cout(s3_345_facout));
full_adder s3_35fa0 ( .A(s1_350_fas), .B(s2_340_facout), .Cin(s2_341_facout), .S(s3_350_fas), .Cout(s3_350_facout));
full_adder s3_35fa1 ( .A(s2_342_facout), .B(s2_343_facout), .Cin(s2_344_facout), .S(s3_351_fas), .Cout(s3_351_facout));
full_adder s3_35fa2 ( .A(s2_345_facout), .B(s2_346_facout), .Cin(s2_347_facout), .S(s3_352_fas), .Cout(s3_352_facout));
full_adder s3_35fa3 ( .A(s2_348_facout), .B(s2_350_fas), .Cin(s2_351_fas), .S(s3_353_fas), .Cout(s3_353_facout));
full_adder s3_35fa4 ( .A(s2_352_fas), .B(s2_353_fas), .Cin(s2_354_fas), .S(s3_354_fas), .Cout(s3_354_facout));
full_adder s3_35fa5 ( .A(s2_355_fas), .B(s2_356_fas), .Cin(s2_357_fas), .S(s3_355_fas), .Cout(s3_355_facout));
full_adder s3_36fa0 ( .A(s1_350_facout), .B(s2_350_facout), .Cin(s2_351_facout), .S(s3_360_fas), .Cout(s3_360_facout));
full_adder s3_36fa1 ( .A(s2_352_facout), .B(s2_353_facout), .Cin(s2_354_facout), .S(s3_361_fas), .Cout(s3_361_facout));
full_adder s3_36fa2 ( .A(s2_355_facout), .B(s2_356_facout), .Cin(s2_357_facout), .S(s3_362_fas), .Cout(s3_362_facout));
full_adder s3_36fa3 ( .A(s2_358_facout), .B(s2_360_fas), .Cin(s2_361_fas), .S(s3_363_fas), .Cout(s3_363_facout));
full_adder s3_36fa4 ( .A(s2_362_fas), .B(s2_363_fas), .Cin(s2_364_fas), .S(s3_364_fas), .Cout(s3_364_facout));
full_adder s3_36fa5 ( .A(s2_365_fas), .B(s2_366_fas), .Cin(s2_367_fas), .S(s3_365_fas), .Cout(s3_365_facout));
full_adder s3_37fa0 ( .A(ps_377), .B(ps_376), .Cin(s2_360_facout), .S(s3_370_fas), .Cout(s3_370_facout));
full_adder s3_37fa1 ( .A(s2_361_facout), .B(s2_362_facout), .Cin(s2_363_facout), .S(s3_371_fas), .Cout(s3_371_facout));
full_adder s3_37fa2 ( .A(s2_364_facout), .B(s2_365_facout), .Cin(s2_366_facout), .S(s3_372_fas), .Cout(s3_372_facout));
full_adder s3_37fa3 ( .A(s2_367_facout), .B(s2_368_facout), .Cin(s2_370_fas), .S(s3_373_fas), .Cout(s3_373_facout));
full_adder s3_37fa4 ( .A(s2_371_fas), .B(s2_372_fas), .Cin(s2_373_fas), .S(s3_374_fas), .Cout(s3_374_facout));
full_adder s3_37fa5 ( .A(s2_374_fas), .B(s2_375_fas), .Cin(s2_376_fas), .S(s3_375_fas), .Cout(s3_375_facout));
full_adder s3_38fa0 ( .A(ps_3810), .B(ps_389), .Cin(ps_388), .S(s3_380_fas), .Cout(s3_380_facout));
full_adder s3_38fa1 ( .A(ps_387), .B(s2_370_facout), .Cin(s2_371_facout), .S(s3_381_fas), .Cout(s3_381_facout));
full_adder s3_38fa2 ( .A(s2_372_facout), .B(s2_373_facout), .Cin(s2_374_facout), .S(s3_382_fas), .Cout(s3_382_facout));
full_adder s3_38fa3 ( .A(s2_375_facout), .B(s2_376_facout), .Cin(s2_377_facout), .S(s3_383_fas), .Cout(s3_383_facout));
full_adder s3_38fa4 ( .A(s2_380_fas), .B(s2_381_fas), .Cin(s2_382_fas), .S(s3_384_fas), .Cout(s3_384_facout));
full_adder s3_38fa5 ( .A(s2_383_fas), .B(s2_384_fas), .Cin(s2_385_fas), .S(s3_385_fas), .Cout(s3_385_facout));
full_adder s3_39fa0 ( .A(ps_3913), .B(ps_3912), .Cin(ps_3911), .S(s3_390_fas), .Cout(s3_390_facout));
full_adder s3_39fa1 ( .A(ps_3910), .B(ps_399), .Cin(ps_398), .S(s3_391_fas), .Cout(s3_391_facout));
full_adder s3_39fa2 ( .A(s2_380_facout), .B(s2_381_facout), .Cin(s2_382_facout), .S(s3_392_fas), .Cout(s3_392_facout));
full_adder s3_39fa3 ( .A(s2_383_facout), .B(s2_384_facout), .Cin(s2_385_facout), .S(s3_393_fas), .Cout(s3_393_facout));
full_adder s3_39fa4 ( .A(s2_386_facout), .B(s2_390_fas), .Cin(s2_391_fas), .S(s3_394_fas), .Cout(s3_394_facout));
full_adder s3_39fa5 ( .A(s2_392_fas), .B(s2_393_fas), .Cin(s2_394_fas), .S(s3_395_fas), .Cout(s3_395_facout));
full_adder s3_40fa0 ( .A(ps_4016), .B(ps_4015), .Cin(ps_4014), .S(s3_400_fas), .Cout(s3_400_facout));
full_adder s3_40fa1 ( .A(ps_4013), .B(ps_4012), .Cin(ps_4011), .S(s3_401_fas), .Cout(s3_401_facout));
full_adder s3_40fa2 ( .A(ps_4010), .B(ps_409), .Cin(s2_390_facout), .S(s3_402_fas), .Cout(s3_402_facout));
full_adder s3_40fa3 ( .A(s2_391_facout), .B(s2_392_facout), .Cin(s2_393_facout), .S(s3_403_fas), .Cout(s3_403_facout));
full_adder s3_40fa4 ( .A(s2_394_facout), .B(s2_395_facout), .Cin(s2_400_fas), .S(s3_404_fas), .Cout(s3_404_facout));
full_adder s3_40fa5 ( .A(s2_401_fas), .B(s2_402_fas), .Cin(s2_403_fas), .S(s3_405_fas), .Cout(s3_405_facout));
full_adder s3_41fa0 ( .A(ps_4119), .B(ps_4118), .Cin(ps_4117), .S(s3_410_fas), .Cout(s3_410_facout));
full_adder s3_41fa1 ( .A(ps_4116), .B(ps_4115), .Cin(ps_4114), .S(s3_411_fas), .Cout(s3_411_facout));
full_adder s3_41fa2 ( .A(ps_4113), .B(ps_4112), .Cin(ps_4111), .S(s3_412_fas), .Cout(s3_412_facout));
full_adder s3_41fa3 ( .A(ps_4110), .B(s2_400_facout), .Cin(s2_401_facout), .S(s3_413_fas), .Cout(s3_413_facout));
full_adder s3_41fa4 ( .A(s2_402_facout), .B(s2_403_facout), .Cin(s2_404_facout), .S(s3_414_fas), .Cout(s3_414_facout));
full_adder s3_41fa5 ( .A(s2_410_fas), .B(s2_411_fas), .Cin(s2_412_fas), .S(s3_415_fas), .Cout(s3_415_facout));
full_adder s3_42fa0 ( .A(ps_4222), .B(ps_4221), .Cin(ps_4220), .S(s3_420_fas), .Cout(s3_420_facout));
full_adder s3_42fa1 ( .A(ps_4219), .B(ps_4218), .Cin(ps_4217), .S(s3_421_fas), .Cout(s3_421_facout));
full_adder s3_42fa2 ( .A(ps_4216), .B(ps_4215), .Cin(ps_4214), .S(s3_422_fas), .Cout(s3_422_facout));
full_adder s3_42fa3 ( .A(ps_4213), .B(ps_4212), .Cin(ps_4211), .S(s3_423_fas), .Cout(s3_423_facout));
full_adder s3_42fa4 ( .A(s2_410_facout), .B(s2_411_facout), .Cin(s2_412_facout), .S(s3_424_fas), .Cout(s3_424_facout));
full_adder s3_42fa5 ( .A(s2_413_facout), .B(s2_420_fas), .Cin(s2_421_fas), .S(s3_425_fas), .Cout(s3_425_facout));
full_adder s3_43fa0 ( .A(ps_4325), .B(ps_4324), .Cin(ps_4323), .S(s3_430_fas), .Cout(s3_430_facout));
full_adder s3_43fa1 ( .A(ps_4322), .B(ps_4321), .Cin(ps_4320), .S(s3_431_fas), .Cout(s3_431_facout));
full_adder s3_43fa2 ( .A(ps_4319), .B(ps_4318), .Cin(ps_4317), .S(s3_432_fas), .Cout(s3_432_facout));
full_adder s3_43fa3 ( .A(ps_4316), .B(ps_4315), .Cin(ps_4314), .S(s3_433_fas), .Cout(s3_433_facout));
full_adder s3_43fa4 ( .A(ps_4313), .B(ps_4312), .Cin(s2_420_facout), .S(s3_434_fas), .Cout(s3_434_facout));
full_adder s3_43fa5 ( .A(s2_421_facout), .B(s2_422_facout), .Cin(s2_430_fas), .S(s3_435_fas), .Cout(s3_435_facout));
full_adder s3_44fa0 ( .A(ps_4428), .B(ps_4427), .Cin(ps_4426), .S(s3_440_fas), .Cout(s3_440_facout));
full_adder s3_44fa1 ( .A(ps_4425), .B(ps_4424), .Cin(ps_4423), .S(s3_441_fas), .Cout(s3_441_facout));
full_adder s3_44fa2 ( .A(ps_4422), .B(ps_4421), .Cin(ps_4420), .S(s3_442_fas), .Cout(s3_442_facout));
full_adder s3_44fa3 ( .A(ps_4419), .B(ps_4418), .Cin(ps_4417), .S(s3_443_fas), .Cout(s3_443_facout));
full_adder s3_44fa4 ( .A(ps_4416), .B(ps_4415), .Cin(ps_4414), .S(s3_444_fas), .Cout(s3_444_facout));
full_adder s3_44fa5 ( .A(ps_4413), .B(s2_430_facout), .Cin(s2_431_facout), .S(s3_445_fas), .Cout(s3_445_facout));
full_adder s3_45fa0 ( .A(ps_4531), .B(ps_4530), .Cin(ps_4529), .S(s3_450_fas), .Cout(s3_450_facout));
full_adder s3_45fa1 ( .A(ps_4528), .B(ps_4527), .Cin(ps_4526), .S(s3_451_fas), .Cout(s3_451_facout));
full_adder s3_45fa2 ( .A(ps_4525), .B(ps_4524), .Cin(ps_4523), .S(s3_452_fas), .Cout(s3_452_facout));
full_adder s3_45fa3 ( .A(ps_4522), .B(ps_4521), .Cin(ps_4520), .S(s3_453_fas), .Cout(s3_453_facout));
full_adder s3_45fa4 ( .A(ps_4519), .B(ps_4518), .Cin(ps_4517), .S(s3_454_fas), .Cout(s3_454_facout));
full_adder s3_45fa5 ( .A(ps_4516), .B(ps_4515), .Cin(ps_4514), .S(s3_455_fas), .Cout(s3_455_facout));
full_adder s3_46fa0 ( .A(ps_4631), .B(ps_4630), .Cin(ps_4629), .S(s3_460_fas), .Cout(s3_460_facout));
full_adder s3_46fa1 ( .A(ps_4628), .B(ps_4627), .Cin(ps_4626), .S(s3_461_fas), .Cout(s3_461_facout));
full_adder s3_46fa2 ( .A(ps_4625), .B(ps_4624), .Cin(ps_4623), .S(s3_462_fas), .Cout(s3_462_facout));
full_adder s3_46fa3 ( .A(ps_4622), .B(ps_4621), .Cin(ps_4620), .S(s3_463_fas), .Cout(s3_463_facout));
full_adder s3_46fa4 ( .A(ps_4619), .B(ps_4618), .Cin(ps_4617), .S(s3_464_fas), .Cout(s3_464_facout));
full_adder s3_47fa0 ( .A(ps_4731), .B(ps_4730), .Cin(ps_4729), .S(s3_470_fas), .Cout(s3_470_facout));
full_adder s3_47fa1 ( .A(ps_4728), .B(ps_4727), .Cin(ps_4726), .S(s3_471_fas), .Cout(s3_471_facout));
full_adder s3_47fa2 ( .A(ps_4725), .B(ps_4724), .Cin(ps_4723), .S(s3_472_fas), .Cout(s3_472_facout));
full_adder s3_47fa3 ( .A(ps_4722), .B(ps_4721), .Cin(ps_4720), .S(s3_473_fas), .Cout(s3_473_facout));
full_adder s3_48fa0 ( .A(ps_4831), .B(ps_4830), .Cin(ps_4829), .S(s3_480_fas), .Cout(s3_480_facout));
full_adder s3_48fa1 ( .A(ps_4828), .B(ps_4827), .Cin(ps_4826), .S(s3_481_fas), .Cout(s3_481_facout));
full_adder s3_48fa2 ( .A(ps_4825), .B(ps_4824), .Cin(ps_4823), .S(s3_482_fas), .Cout(s3_482_facout));
full_adder s3_49fa0 ( .A(ps_4931), .B(ps_4930), .Cin(ps_4929), .S(s3_490_fas), .Cout(s3_490_facout));
full_adder s3_49fa1 ( .A(ps_4928), .B(ps_4927), .Cin(ps_4926), .S(s3_491_fas), .Cout(s3_491_facout));
full_adder s3_50fa0 ( .A(ps_5031), .B(ps_5030), .Cin(ps_5029), .S(s3_500_fas), .Cout(s3_500_facout));
logic s4_90_hacout, s4_90_has, s4_100_facout, s4_100_fas, s4_100_hacout, s4_100_has, s4_110_facout, s4_110_fas, s4_111_facout, s4_111_fas, s4_110_hacout, s4_110_has, s4_120_facout, s4_120_fas, s4_121_facout, s4_121_fas, s4_122_facout, s4_122_fas, s4_120_hacout, s4_120_has, s4_130_facout, s4_130_fas, s4_131_facout, s4_131_fas, s4_132_facout, s4_132_fas, s4_133_facout, s4_133_fas, s4_140_facout, s4_140_fas, s4_141_facout, s4_141_fas, s4_142_facout, s4_142_fas, s4_143_facout, s4_143_fas, s4_150_facout, s4_150_fas, s4_151_facout, s4_151_fas, s4_152_facout, s4_152_fas, s4_153_facout, s4_153_fas, s4_160_facout, s4_160_fas, s4_161_facout, s4_161_fas, s4_162_facout, s4_162_fas, s4_163_facout, s4_163_fas, s4_170_facout, s4_170_fas, s4_171_facout, s4_171_fas, s4_172_facout, s4_172_fas, s4_173_facout, s4_173_fas, s4_180_facout, s4_180_fas, s4_181_facout, s4_181_fas, s4_182_facout, s4_182_fas, s4_183_facout, s4_183_fas, s4_190_facout, s4_190_fas, s4_191_facout, s4_191_fas, s4_192_facout, s4_192_fas, s4_193_facout, s4_193_fas, s4_200_facout, s4_200_fas, s4_201_facout, s4_201_fas, s4_202_facout, s4_202_fas, s4_203_facout, s4_203_fas, s4_210_facout, s4_210_fas, s4_211_facout, s4_211_fas, s4_212_facout, s4_212_fas, s4_213_facout, s4_213_fas, s4_220_facout, s4_220_fas, s4_221_facout, s4_221_fas, s4_222_facout, s4_222_fas, s4_223_facout, s4_223_fas, s4_230_facout, s4_230_fas, s4_231_facout, s4_231_fas, s4_232_facout, s4_232_fas, s4_233_facout, s4_233_fas, s4_240_facout, s4_240_fas, s4_241_facout, s4_241_fas, s4_242_facout, s4_242_fas, s4_243_facout, s4_243_fas, s4_250_facout, s4_250_fas, s4_251_facout, s4_251_fas, s4_252_facout, s4_252_fas, s4_253_facout, s4_253_fas, s4_260_facout, s4_260_fas, s4_261_facout, s4_261_fas, s4_262_facout, s4_262_fas, s4_263_facout, s4_263_fas, s4_270_facout, s4_270_fas, s4_271_facout, s4_271_fas, s4_272_facout, s4_272_fas, s4_273_facout, s4_273_fas, s4_280_facout, s4_280_fas, s4_281_facout, s4_281_fas, s4_282_facout, s4_282_fas, s4_283_facout, s4_283_fas, s4_290_facout, s4_290_fas, s4_291_facout, s4_291_fas, s4_292_facout, s4_292_fas, s4_293_facout, s4_293_fas, s4_300_facout, s4_300_fas, s4_301_facout, s4_301_fas, s4_302_facout, s4_302_fas, s4_303_facout, s4_303_fas, s4_310_facout, s4_310_fas, s4_311_facout, s4_311_fas, s4_312_facout, s4_312_fas, s4_313_facout, s4_313_fas, s4_320_facout, s4_320_fas, s4_321_facout, s4_321_fas, s4_322_facout, s4_322_fas, s4_323_facout, s4_323_fas, s4_330_facout, s4_330_fas, s4_331_facout, s4_331_fas, s4_332_facout, s4_332_fas, s4_333_facout, s4_333_fas, s4_340_facout, s4_340_fas, s4_341_facout, s4_341_fas, s4_342_facout, s4_342_fas, s4_343_facout, s4_343_fas, s4_350_facout, s4_350_fas, s4_351_facout, s4_351_fas, s4_352_facout, s4_352_fas, s4_353_facout, s4_353_fas, s4_360_facout, s4_360_fas, s4_361_facout, s4_361_fas, s4_362_facout, s4_362_fas, s4_363_facout, s4_363_fas, s4_370_facout, s4_370_fas, s4_371_facout, s4_371_fas, s4_372_facout, s4_372_fas, s4_373_facout, s4_373_fas, s4_380_facout, s4_380_fas, s4_381_facout, s4_381_fas, s4_382_facout, s4_382_fas, s4_383_facout, s4_383_fas, s4_390_facout, s4_390_fas, s4_391_facout, s4_391_fas, s4_392_facout, s4_392_fas, s4_393_facout, s4_393_fas, s4_400_facout, s4_400_fas, s4_401_facout, s4_401_fas, s4_402_facout, s4_402_fas, s4_403_facout, s4_403_fas, s4_410_facout, s4_410_fas, s4_411_facout, s4_411_fas, s4_412_facout, s4_412_fas, s4_413_facout, s4_413_fas, s4_420_facout, s4_420_fas, s4_421_facout, s4_421_fas, s4_422_facout, s4_422_fas, s4_423_facout, s4_423_fas, s4_430_facout, s4_430_fas, s4_431_facout, s4_431_fas, s4_432_facout, s4_432_fas, s4_433_facout, s4_433_fas, s4_440_facout, s4_440_fas, s4_441_facout, s4_441_fas, s4_442_facout, s4_442_fas, s4_443_facout, s4_443_fas, s4_450_facout, s4_450_fas, s4_451_facout, s4_451_fas, s4_452_facout, s4_452_fas, s4_453_facout, s4_453_fas, s4_460_facout, s4_460_fas, s4_461_facout, s4_461_fas, s4_462_facout, s4_462_fas, s4_463_facout, s4_463_fas, s4_470_facout, s4_470_fas, s4_471_facout, s4_471_fas, s4_472_facout, s4_472_fas, s4_473_facout, s4_473_fas, s4_480_facout, s4_480_fas, s4_481_facout, s4_481_fas, s4_482_facout, s4_482_fas, s4_483_facout, s4_483_fas, s4_490_facout, s4_490_fas, s4_491_facout, s4_491_fas, s4_492_facout, s4_492_fas, s4_493_facout, s4_493_fas, s4_500_facout, s4_500_fas, s4_501_facout, s4_501_fas, s4_502_facout, s4_502_fas, s4_503_facout, s4_503_fas, s4_510_facout, s4_510_fas, s4_511_facout, s4_511_fas, s4_512_facout, s4_512_fas, s4_513_facout, s4_513_fas, s4_520_facout, s4_520_fas, s4_521_facout, s4_521_fas, s4_522_facout, s4_522_fas, s4_530_facout, s4_530_fas, s4_531_facout, s4_531_fas, s4_540_facout, s4_540_fas;
/* ========================= Stage 4 ========================= */
half_adder s4_9ha0 ( .A(ps_99), .B(ps_98), .S(s4_90_has), .Cout(s4_90_hacout));
full_adder s4_10fa0 ( .A(ps_1010), .B(ps_109), .Cin(ps_108), .S(s4_100_fas), .Cout(s4_100_facout));
half_adder s4_10ha0 ( .A(ps_107), .B(ps_106), .S(s4_100_has), .Cout(s4_100_hacout));
full_adder s4_11fa0 ( .A(ps_1111), .B(ps_1110), .Cin(ps_119), .S(s4_110_fas), .Cout(s4_110_facout));
full_adder s4_11fa1 ( .A(ps_118), .B(ps_117), .Cin(ps_116), .S(s4_111_fas), .Cout(s4_111_facout));
half_adder s4_11ha0 ( .A(ps_115), .B(ps_114), .S(s4_110_has), .Cout(s4_110_hacout));
full_adder s4_12fa0 ( .A(ps_1212), .B(ps_1211), .Cin(ps_1210), .S(s4_120_fas), .Cout(s4_120_facout));
full_adder s4_12fa1 ( .A(ps_129), .B(ps_128), .Cin(ps_127), .S(s4_121_fas), .Cout(s4_121_facout));
full_adder s4_12fa2 ( .A(ps_126), .B(ps_125), .Cin(ps_124), .S(s4_122_fas), .Cout(s4_122_facout));
half_adder s4_12ha0 ( .A(ps_123), .B(ps_122), .S(s4_120_has), .Cout(s4_120_hacout));
full_adder s4_13fa0 ( .A(ps_1311), .B(ps_1310), .Cin(ps_139), .S(s4_130_fas), .Cout(s4_130_facout));
full_adder s4_13fa1 ( .A(ps_138), .B(ps_137), .Cin(ps_136), .S(s4_131_fas), .Cout(s4_131_facout));
full_adder s4_13fa2 ( .A(ps_135), .B(ps_134), .Cin(ps_133), .S(s4_132_fas), .Cout(s4_132_facout));
full_adder s4_13fa3 ( .A(ps_132), .B(ps_131), .Cin(ps_130), .S(s4_133_fas), .Cout(s4_133_facout));
full_adder s4_14fa0 ( .A(ps_149), .B(ps_148), .Cin(ps_147), .S(s4_140_fas), .Cout(s4_140_facout));
full_adder s4_14fa1 ( .A(ps_146), .B(ps_145), .Cin(ps_144), .S(s4_141_fas), .Cout(s4_141_facout));
full_adder s4_14fa2 ( .A(ps_143), .B(ps_142), .Cin(ps_141), .S(s4_142_fas), .Cout(s4_142_facout));
full_adder s4_14fa3 ( .A(ps_140), .B(s3_130_hacout), .Cin(s3_140_fas), .S(s4_143_fas), .Cout(s4_143_facout));
full_adder s4_15fa0 ( .A(ps_157), .B(ps_156), .Cin(ps_155), .S(s4_150_fas), .Cout(s4_150_facout));
full_adder s4_15fa1 ( .A(ps_154), .B(ps_153), .Cin(ps_152), .S(s4_151_fas), .Cout(s4_151_facout));
full_adder s4_15fa2 ( .A(ps_151), .B(ps_150), .Cin(s3_140_facout), .S(s4_152_fas), .Cout(s4_152_facout));
full_adder s4_15fa3 ( .A(s3_140_hacout), .B(s3_150_fas), .Cin(s3_151_fas), .S(s4_153_fas), .Cout(s4_153_facout));
full_adder s4_16fa0 ( .A(ps_165), .B(ps_164), .Cin(ps_163), .S(s4_160_fas), .Cout(s4_160_facout));
full_adder s4_16fa1 ( .A(ps_162), .B(ps_161), .Cin(ps_160), .S(s4_161_fas), .Cout(s4_161_facout));
full_adder s4_16fa2 ( .A(s3_150_facout), .B(s3_151_facout), .Cin(s3_150_hacout), .S(s4_162_fas), .Cout(s4_162_facout));
full_adder s4_16fa3 ( .A(s3_160_fas), .B(s3_161_fas), .Cin(s3_162_fas), .S(s4_163_fas), .Cout(s4_163_facout));
full_adder s4_17fa0 ( .A(ps_173), .B(ps_172), .Cin(ps_171), .S(s4_170_fas), .Cout(s4_170_facout));
full_adder s4_17fa1 ( .A(ps_170), .B(s3_160_facout), .Cin(s3_161_facout), .S(s4_171_fas), .Cout(s4_171_facout));
full_adder s4_17fa2 ( .A(s3_162_facout), .B(s3_160_hacout), .Cin(s3_170_fas), .S(s4_172_fas), .Cout(s4_172_facout));
full_adder s4_17fa3 ( .A(s3_171_fas), .B(s3_172_fas), .Cin(s3_173_fas), .S(s4_173_fas), .Cout(s4_173_facout));
full_adder s4_18fa0 ( .A(ps_181), .B(ps_180), .Cin(s3_170_facout), .S(s4_180_fas), .Cout(s4_180_facout));
full_adder s4_18fa1 ( .A(s3_171_facout), .B(s3_172_facout), .Cin(s3_173_facout), .S(s4_181_fas), .Cout(s4_181_facout));
full_adder s4_18fa2 ( .A(s3_170_hacout), .B(s3_180_fas), .Cin(s3_181_fas), .S(s4_182_fas), .Cout(s4_182_facout));
full_adder s4_18fa3 ( .A(s3_182_fas), .B(s3_183_fas), .Cin(s3_184_fas), .S(s4_183_fas), .Cout(s4_183_facout));
full_adder s4_19fa0 ( .A(s2_190_has), .B(s3_180_facout), .Cin(s3_181_facout), .S(s4_190_fas), .Cout(s4_190_facout));
full_adder s4_19fa1 ( .A(s3_182_facout), .B(s3_183_facout), .Cin(s3_184_facout), .S(s4_191_fas), .Cout(s4_191_facout));
full_adder s4_19fa2 ( .A(s3_180_hacout), .B(s3_190_fas), .Cin(s3_191_fas), .S(s4_192_fas), .Cout(s4_192_facout));
full_adder s4_19fa3 ( .A(s3_192_fas), .B(s3_193_fas), .Cin(s3_194_fas), .S(s4_193_fas), .Cout(s4_193_facout));
full_adder s4_20fa0 ( .A(s2_200_has), .B(s3_190_facout), .Cin(s3_191_facout), .S(s4_200_fas), .Cout(s4_200_facout));
full_adder s4_20fa1 ( .A(s3_192_facout), .B(s3_193_facout), .Cin(s3_194_facout), .S(s4_201_fas), .Cout(s4_201_facout));
full_adder s4_20fa2 ( .A(s3_195_facout), .B(s3_200_fas), .Cin(s3_201_fas), .S(s4_202_fas), .Cout(s4_202_facout));
full_adder s4_20fa3 ( .A(s3_202_fas), .B(s3_203_fas), .Cin(s3_204_fas), .S(s4_203_fas), .Cout(s4_203_facout));
full_adder s4_21fa0 ( .A(s2_210_has), .B(s3_200_facout), .Cin(s3_201_facout), .S(s4_210_fas), .Cout(s4_210_facout));
full_adder s4_21fa1 ( .A(s3_202_facout), .B(s3_203_facout), .Cin(s3_204_facout), .S(s4_211_fas), .Cout(s4_211_facout));
full_adder s4_21fa2 ( .A(s3_205_facout), .B(s3_210_fas), .Cin(s3_211_fas), .S(s4_212_fas), .Cout(s4_212_facout));
full_adder s4_21fa3 ( .A(s3_212_fas), .B(s3_213_fas), .Cin(s3_214_fas), .S(s4_213_fas), .Cout(s4_213_facout));
full_adder s4_22fa0 ( .A(s2_220_has), .B(s3_210_facout), .Cin(s3_211_facout), .S(s4_220_fas), .Cout(s4_220_facout));
full_adder s4_22fa1 ( .A(s3_212_facout), .B(s3_213_facout), .Cin(s3_214_facout), .S(s4_221_fas), .Cout(s4_221_facout));
full_adder s4_22fa2 ( .A(s3_215_facout), .B(s3_220_fas), .Cin(s3_221_fas), .S(s4_222_fas), .Cout(s4_222_facout));
full_adder s4_22fa3 ( .A(s3_222_fas), .B(s3_223_fas), .Cin(s3_224_fas), .S(s4_223_fas), .Cout(s4_223_facout));
full_adder s4_23fa0 ( .A(s2_230_has), .B(s3_220_facout), .Cin(s3_221_facout), .S(s4_230_fas), .Cout(s4_230_facout));
full_adder s4_23fa1 ( .A(s3_222_facout), .B(s3_223_facout), .Cin(s3_224_facout), .S(s4_231_fas), .Cout(s4_231_facout));
full_adder s4_23fa2 ( .A(s3_225_facout), .B(s3_230_fas), .Cin(s3_231_fas), .S(s4_232_fas), .Cout(s4_232_facout));
full_adder s4_23fa3 ( .A(s3_232_fas), .B(s3_233_fas), .Cin(s3_234_fas), .S(s4_233_fas), .Cout(s4_233_facout));
full_adder s4_24fa0 ( .A(s2_240_has), .B(s3_230_facout), .Cin(s3_231_facout), .S(s4_240_fas), .Cout(s4_240_facout));
full_adder s4_24fa1 ( .A(s3_232_facout), .B(s3_233_facout), .Cin(s3_234_facout), .S(s4_241_fas), .Cout(s4_241_facout));
full_adder s4_24fa2 ( .A(s3_235_facout), .B(s3_240_fas), .Cin(s3_241_fas), .S(s4_242_fas), .Cout(s4_242_facout));
full_adder s4_24fa3 ( .A(s3_242_fas), .B(s3_243_fas), .Cin(s3_244_fas), .S(s4_243_fas), .Cout(s4_243_facout));
full_adder s4_25fa0 ( .A(s2_250_has), .B(s3_240_facout), .Cin(s3_241_facout), .S(s4_250_fas), .Cout(s4_250_facout));
full_adder s4_25fa1 ( .A(s3_242_facout), .B(s3_243_facout), .Cin(s3_244_facout), .S(s4_251_fas), .Cout(s4_251_facout));
full_adder s4_25fa2 ( .A(s3_245_facout), .B(s3_250_fas), .Cin(s3_251_fas), .S(s4_252_fas), .Cout(s4_252_facout));
full_adder s4_25fa3 ( .A(s3_252_fas), .B(s3_253_fas), .Cin(s3_254_fas), .S(s4_253_fas), .Cout(s4_253_facout));
full_adder s4_26fa0 ( .A(s2_260_has), .B(s3_250_facout), .Cin(s3_251_facout), .S(s4_260_fas), .Cout(s4_260_facout));
full_adder s4_26fa1 ( .A(s3_252_facout), .B(s3_253_facout), .Cin(s3_254_facout), .S(s4_261_fas), .Cout(s4_261_facout));
full_adder s4_26fa2 ( .A(s3_255_facout), .B(s3_260_fas), .Cin(s3_261_fas), .S(s4_262_fas), .Cout(s4_262_facout));
full_adder s4_26fa3 ( .A(s3_262_fas), .B(s3_263_fas), .Cin(s3_264_fas), .S(s4_263_fas), .Cout(s4_263_facout));
full_adder s4_27fa0 ( .A(s2_270_has), .B(s3_260_facout), .Cin(s3_261_facout), .S(s4_270_fas), .Cout(s4_270_facout));
full_adder s4_27fa1 ( .A(s3_262_facout), .B(s3_263_facout), .Cin(s3_264_facout), .S(s4_271_fas), .Cout(s4_271_facout));
full_adder s4_27fa2 ( .A(s3_265_facout), .B(s3_270_fas), .Cin(s3_271_fas), .S(s4_272_fas), .Cout(s4_272_facout));
full_adder s4_27fa3 ( .A(s3_272_fas), .B(s3_273_fas), .Cin(s3_274_fas), .S(s4_273_fas), .Cout(s4_273_facout));
full_adder s4_28fa0 ( .A(s2_288_fas), .B(s3_270_facout), .Cin(s3_271_facout), .S(s4_280_fas), .Cout(s4_280_facout));
full_adder s4_28fa1 ( .A(s3_272_facout), .B(s3_273_facout), .Cin(s3_274_facout), .S(s4_281_fas), .Cout(s4_281_facout));
full_adder s4_28fa2 ( .A(s3_275_facout), .B(s3_280_fas), .Cin(s3_281_fas), .S(s4_282_fas), .Cout(s4_282_facout));
full_adder s4_28fa3 ( .A(s3_282_fas), .B(s3_283_fas), .Cin(s3_284_fas), .S(s4_283_fas), .Cout(s4_283_facout));
full_adder s4_29fa0 ( .A(s2_298_fas), .B(s3_280_facout), .Cin(s3_281_facout), .S(s4_290_fas), .Cout(s4_290_facout));
full_adder s4_29fa1 ( .A(s3_282_facout), .B(s3_283_facout), .Cin(s3_284_facout), .S(s4_291_fas), .Cout(s4_291_facout));
full_adder s4_29fa2 ( .A(s3_285_facout), .B(s3_290_fas), .Cin(s3_291_fas), .S(s4_292_fas), .Cout(s4_292_facout));
full_adder s4_29fa3 ( .A(s3_292_fas), .B(s3_293_fas), .Cin(s3_294_fas), .S(s4_293_fas), .Cout(s4_293_facout));
full_adder s4_30fa0 ( .A(s2_308_fas), .B(s3_290_facout), .Cin(s3_291_facout), .S(s4_300_fas), .Cout(s4_300_facout));
full_adder s4_30fa1 ( .A(s3_292_facout), .B(s3_293_facout), .Cin(s3_294_facout), .S(s4_301_fas), .Cout(s4_301_facout));
full_adder s4_30fa2 ( .A(s3_295_facout), .B(s3_300_fas), .Cin(s3_301_fas), .S(s4_302_fas), .Cout(s4_302_facout));
full_adder s4_30fa3 ( .A(s3_302_fas), .B(s3_303_fas), .Cin(s3_304_fas), .S(s4_303_fas), .Cout(s4_303_facout));
full_adder s4_31fa0 ( .A(s2_318_fas), .B(s3_300_facout), .Cin(s3_301_facout), .S(s4_310_fas), .Cout(s4_310_facout));
full_adder s4_31fa1 ( .A(s3_302_facout), .B(s3_303_facout), .Cin(s3_304_facout), .S(s4_311_fas), .Cout(s4_311_facout));
full_adder s4_31fa2 ( .A(s3_305_facout), .B(s3_310_fas), .Cin(s3_311_fas), .S(s4_312_fas), .Cout(s4_312_facout));
full_adder s4_31fa3 ( .A(s3_312_fas), .B(s3_313_fas), .Cin(s3_314_fas), .S(s4_313_fas), .Cout(s4_313_facout));
full_adder s4_32fa0 ( .A(s2_328_fas), .B(s3_310_facout), .Cin(s3_311_facout), .S(s4_320_fas), .Cout(s4_320_facout));
full_adder s4_32fa1 ( .A(s3_312_facout), .B(s3_313_facout), .Cin(s3_314_facout), .S(s4_321_fas), .Cout(s4_321_facout));
full_adder s4_32fa2 ( .A(s3_315_facout), .B(s3_320_fas), .Cin(s3_321_fas), .S(s4_322_fas), .Cout(s4_322_facout));
full_adder s4_32fa3 ( .A(s3_322_fas), .B(s3_323_fas), .Cin(s3_324_fas), .S(s4_323_fas), .Cout(s4_323_facout));
full_adder s4_33fa0 ( .A(s2_338_fas), .B(s3_320_facout), .Cin(s3_321_facout), .S(s4_330_fas), .Cout(s4_330_facout));
full_adder s4_33fa1 ( .A(s3_322_facout), .B(s3_323_facout), .Cin(s3_324_facout), .S(s4_331_fas), .Cout(s4_331_facout));
full_adder s4_33fa2 ( .A(s3_325_facout), .B(s3_330_fas), .Cin(s3_331_fas), .S(s4_332_fas), .Cout(s4_332_facout));
full_adder s4_33fa3 ( .A(s3_332_fas), .B(s3_333_fas), .Cin(s3_334_fas), .S(s4_333_fas), .Cout(s4_333_facout));
full_adder s4_34fa0 ( .A(s2_348_fas), .B(s3_330_facout), .Cin(s3_331_facout), .S(s4_340_fas), .Cout(s4_340_facout));
full_adder s4_34fa1 ( .A(s3_332_facout), .B(s3_333_facout), .Cin(s3_334_facout), .S(s4_341_fas), .Cout(s4_341_facout));
full_adder s4_34fa2 ( .A(s3_335_facout), .B(s3_340_fas), .Cin(s3_341_fas), .S(s4_342_fas), .Cout(s4_342_facout));
full_adder s4_34fa3 ( .A(s3_342_fas), .B(s3_343_fas), .Cin(s3_344_fas), .S(s4_343_fas), .Cout(s4_343_facout));
full_adder s4_35fa0 ( .A(s2_358_fas), .B(s3_340_facout), .Cin(s3_341_facout), .S(s4_350_fas), .Cout(s4_350_facout));
full_adder s4_35fa1 ( .A(s3_342_facout), .B(s3_343_facout), .Cin(s3_344_facout), .S(s4_351_fas), .Cout(s4_351_facout));
full_adder s4_35fa2 ( .A(s3_345_facout), .B(s3_350_fas), .Cin(s3_351_fas), .S(s4_352_fas), .Cout(s4_352_facout));
full_adder s4_35fa3 ( .A(s3_352_fas), .B(s3_353_fas), .Cin(s3_354_fas), .S(s4_353_fas), .Cout(s4_353_facout));
full_adder s4_36fa0 ( .A(s2_368_fas), .B(s3_350_facout), .Cin(s3_351_facout), .S(s4_360_fas), .Cout(s4_360_facout));
full_adder s4_36fa1 ( .A(s3_352_facout), .B(s3_353_facout), .Cin(s3_354_facout), .S(s4_361_fas), .Cout(s4_361_facout));
full_adder s4_36fa2 ( .A(s3_355_facout), .B(s3_360_fas), .Cin(s3_361_fas), .S(s4_362_fas), .Cout(s4_362_facout));
full_adder s4_36fa3 ( .A(s3_362_fas), .B(s3_363_fas), .Cin(s3_364_fas), .S(s4_363_fas), .Cout(s4_363_facout));
full_adder s4_37fa0 ( .A(s2_377_fas), .B(s3_360_facout), .Cin(s3_361_facout), .S(s4_370_fas), .Cout(s4_370_facout));
full_adder s4_37fa1 ( .A(s3_362_facout), .B(s3_363_facout), .Cin(s3_364_facout), .S(s4_371_fas), .Cout(s4_371_facout));
full_adder s4_37fa2 ( .A(s3_365_facout), .B(s3_370_fas), .Cin(s3_371_fas), .S(s4_372_fas), .Cout(s4_372_facout));
full_adder s4_37fa3 ( .A(s3_372_fas), .B(s3_373_fas), .Cin(s3_374_fas), .S(s4_373_fas), .Cout(s4_373_facout));
full_adder s4_38fa0 ( .A(s2_386_fas), .B(s3_370_facout), .Cin(s3_371_facout), .S(s4_380_fas), .Cout(s4_380_facout));
full_adder s4_38fa1 ( .A(s3_372_facout), .B(s3_373_facout), .Cin(s3_374_facout), .S(s4_381_fas), .Cout(s4_381_facout));
full_adder s4_38fa2 ( .A(s3_375_facout), .B(s3_380_fas), .Cin(s3_381_fas), .S(s4_382_fas), .Cout(s4_382_facout));
full_adder s4_38fa3 ( .A(s3_382_fas), .B(s3_383_fas), .Cin(s3_384_fas), .S(s4_383_fas), .Cout(s4_383_facout));
full_adder s4_39fa0 ( .A(s2_395_fas), .B(s3_380_facout), .Cin(s3_381_facout), .S(s4_390_fas), .Cout(s4_390_facout));
full_adder s4_39fa1 ( .A(s3_382_facout), .B(s3_383_facout), .Cin(s3_384_facout), .S(s4_391_fas), .Cout(s4_391_facout));
full_adder s4_39fa2 ( .A(s3_385_facout), .B(s3_390_fas), .Cin(s3_391_fas), .S(s4_392_fas), .Cout(s4_392_facout));
full_adder s4_39fa3 ( .A(s3_392_fas), .B(s3_393_fas), .Cin(s3_394_fas), .S(s4_393_fas), .Cout(s4_393_facout));
full_adder s4_40fa0 ( .A(s2_404_fas), .B(s3_390_facout), .Cin(s3_391_facout), .S(s4_400_fas), .Cout(s4_400_facout));
full_adder s4_40fa1 ( .A(s3_392_facout), .B(s3_393_facout), .Cin(s3_394_facout), .S(s4_401_fas), .Cout(s4_401_facout));
full_adder s4_40fa2 ( .A(s3_395_facout), .B(s3_400_fas), .Cin(s3_401_fas), .S(s4_402_fas), .Cout(s4_402_facout));
full_adder s4_40fa3 ( .A(s3_402_fas), .B(s3_403_fas), .Cin(s3_404_fas), .S(s4_403_fas), .Cout(s4_403_facout));
full_adder s4_41fa0 ( .A(s2_413_fas), .B(s3_400_facout), .Cin(s3_401_facout), .S(s4_410_fas), .Cout(s4_410_facout));
full_adder s4_41fa1 ( .A(s3_402_facout), .B(s3_403_facout), .Cin(s3_404_facout), .S(s4_411_fas), .Cout(s4_411_facout));
full_adder s4_41fa2 ( .A(s3_405_facout), .B(s3_410_fas), .Cin(s3_411_fas), .S(s4_412_fas), .Cout(s4_412_facout));
full_adder s4_41fa3 ( .A(s3_412_fas), .B(s3_413_fas), .Cin(s3_414_fas), .S(s4_413_fas), .Cout(s4_413_facout));
full_adder s4_42fa0 ( .A(s2_422_fas), .B(s3_410_facout), .Cin(s3_411_facout), .S(s4_420_fas), .Cout(s4_420_facout));
full_adder s4_42fa1 ( .A(s3_412_facout), .B(s3_413_facout), .Cin(s3_414_facout), .S(s4_421_fas), .Cout(s4_421_facout));
full_adder s4_42fa2 ( .A(s3_415_facout), .B(s3_420_fas), .Cin(s3_421_fas), .S(s4_422_fas), .Cout(s4_422_facout));
full_adder s4_42fa3 ( .A(s3_422_fas), .B(s3_423_fas), .Cin(s3_424_fas), .S(s4_423_fas), .Cout(s4_423_facout));
full_adder s4_43fa0 ( .A(s2_431_fas), .B(s3_420_facout), .Cin(s3_421_facout), .S(s4_430_fas), .Cout(s4_430_facout));
full_adder s4_43fa1 ( .A(s3_422_facout), .B(s3_423_facout), .Cin(s3_424_facout), .S(s4_431_fas), .Cout(s4_431_facout));
full_adder s4_43fa2 ( .A(s3_425_facout), .B(s3_430_fas), .Cin(s3_431_fas), .S(s4_432_fas), .Cout(s4_432_facout));
full_adder s4_43fa3 ( .A(s3_432_fas), .B(s3_433_fas), .Cin(s3_434_fas), .S(s4_433_fas), .Cout(s4_433_facout));
full_adder s4_44fa0 ( .A(s2_440_fas), .B(s3_430_facout), .Cin(s3_431_facout), .S(s4_440_fas), .Cout(s4_440_facout));
full_adder s4_44fa1 ( .A(s3_432_facout), .B(s3_433_facout), .Cin(s3_434_facout), .S(s4_441_fas), .Cout(s4_441_facout));
full_adder s4_44fa2 ( .A(s3_435_facout), .B(s3_440_fas), .Cin(s3_441_fas), .S(s4_442_fas), .Cout(s4_442_facout));
full_adder s4_44fa3 ( .A(s3_442_fas), .B(s3_443_fas), .Cin(s3_444_fas), .S(s4_443_fas), .Cout(s4_443_facout));
full_adder s4_45fa0 ( .A(s2_440_facout), .B(s3_440_facout), .Cin(s3_441_facout), .S(s4_450_fas), .Cout(s4_450_facout));
full_adder s4_45fa1 ( .A(s3_442_facout), .B(s3_443_facout), .Cin(s3_444_facout), .S(s4_451_fas), .Cout(s4_451_facout));
full_adder s4_45fa2 ( .A(s3_445_facout), .B(s3_450_fas), .Cin(s3_451_fas), .S(s4_452_fas), .Cout(s4_452_facout));
full_adder s4_45fa3 ( .A(s3_452_fas), .B(s3_453_fas), .Cin(s3_454_fas), .S(s4_453_fas), .Cout(s4_453_facout));
full_adder s4_46fa0 ( .A(ps_4616), .B(ps_4615), .Cin(s3_450_facout), .S(s4_460_fas), .Cout(s4_460_facout));
full_adder s4_46fa1 ( .A(s3_451_facout), .B(s3_452_facout), .Cin(s3_453_facout), .S(s4_461_fas), .Cout(s4_461_facout));
full_adder s4_46fa2 ( .A(s3_454_facout), .B(s3_455_facout), .Cin(s3_460_fas), .S(s4_462_fas), .Cout(s4_462_facout));
full_adder s4_46fa3 ( .A(s3_461_fas), .B(s3_462_fas), .Cin(s3_463_fas), .S(s4_463_fas), .Cout(s4_463_facout));
full_adder s4_47fa0 ( .A(ps_4719), .B(ps_4718), .Cin(ps_4717), .S(s4_470_fas), .Cout(s4_470_facout));
full_adder s4_47fa1 ( .A(ps_4716), .B(s3_460_facout), .Cin(s3_461_facout), .S(s4_471_fas), .Cout(s4_471_facout));
full_adder s4_47fa2 ( .A(s3_462_facout), .B(s3_463_facout), .Cin(s3_464_facout), .S(s4_472_fas), .Cout(s4_472_facout));
full_adder s4_47fa3 ( .A(s3_470_fas), .B(s3_471_fas), .Cin(s3_472_fas), .S(s4_473_fas), .Cout(s4_473_facout));
full_adder s4_48fa0 ( .A(ps_4822), .B(ps_4821), .Cin(ps_4820), .S(s4_480_fas), .Cout(s4_480_facout));
full_adder s4_48fa1 ( .A(ps_4819), .B(ps_4818), .Cin(ps_4817), .S(s4_481_fas), .Cout(s4_481_facout));
full_adder s4_48fa2 ( .A(s3_470_facout), .B(s3_471_facout), .Cin(s3_472_facout), .S(s4_482_fas), .Cout(s4_482_facout));
full_adder s4_48fa3 ( .A(s3_473_facout), .B(s3_480_fas), .Cin(s3_481_fas), .S(s4_483_fas), .Cout(s4_483_facout));
full_adder s4_49fa0 ( .A(ps_4925), .B(ps_4924), .Cin(ps_4923), .S(s4_490_fas), .Cout(s4_490_facout));
full_adder s4_49fa1 ( .A(ps_4922), .B(ps_4921), .Cin(ps_4920), .S(s4_491_fas), .Cout(s4_491_facout));
full_adder s4_49fa2 ( .A(ps_4919), .B(ps_4918), .Cin(s3_480_facout), .S(s4_492_fas), .Cout(s4_492_facout));
full_adder s4_49fa3 ( .A(s3_481_facout), .B(s3_482_facout), .Cin(s3_490_fas), .S(s4_493_fas), .Cout(s4_493_facout));
full_adder s4_50fa0 ( .A(ps_5028), .B(ps_5027), .Cin(ps_5026), .S(s4_500_fas), .Cout(s4_500_facout));
full_adder s4_50fa1 ( .A(ps_5025), .B(ps_5024), .Cin(ps_5023), .S(s4_501_fas), .Cout(s4_501_facout));
full_adder s4_50fa2 ( .A(ps_5022), .B(ps_5021), .Cin(ps_5020), .S(s4_502_fas), .Cout(s4_502_facout));
full_adder s4_50fa3 ( .A(ps_5019), .B(s3_490_facout), .Cin(s3_491_facout), .S(s4_503_fas), .Cout(s4_503_facout));
full_adder s4_51fa0 ( .A(ps_5131), .B(ps_5130), .Cin(ps_5129), .S(s4_510_fas), .Cout(s4_510_facout));
full_adder s4_51fa1 ( .A(ps_5128), .B(ps_5127), .Cin(ps_5126), .S(s4_511_fas), .Cout(s4_511_facout));
full_adder s4_51fa2 ( .A(ps_5125), .B(ps_5124), .Cin(ps_5123), .S(s4_512_fas), .Cout(s4_512_facout));
full_adder s4_51fa3 ( .A(ps_5122), .B(ps_5121), .Cin(ps_5120), .S(s4_513_fas), .Cout(s4_513_facout));
full_adder s4_52fa0 ( .A(ps_5231), .B(ps_5230), .Cin(ps_5229), .S(s4_520_fas), .Cout(s4_520_facout));
full_adder s4_52fa1 ( .A(ps_5228), .B(ps_5227), .Cin(ps_5226), .S(s4_521_fas), .Cout(s4_521_facout));
full_adder s4_52fa2 ( .A(ps_5225), .B(ps_5224), .Cin(ps_5223), .S(s4_522_fas), .Cout(s4_522_facout));
full_adder s4_53fa0 ( .A(ps_5331), .B(ps_5330), .Cin(ps_5329), .S(s4_530_fas), .Cout(s4_530_facout));
full_adder s4_53fa1 ( .A(ps_5328), .B(ps_5327), .Cin(ps_5326), .S(s4_531_fas), .Cout(s4_531_facout));
full_adder s4_54fa0 ( .A(ps_5431), .B(ps_5430), .Cin(ps_5429), .S(s4_540_fas), .Cout(s4_540_facout));
logic s5_60_hacout, s5_60_has, s5_70_facout, s5_70_fas, s5_70_hacout, s5_70_has, s5_80_facout, s5_80_fas, s5_81_facout, s5_81_fas, s5_80_hacout, s5_80_has, s5_90_facout, s5_90_fas, s5_91_facout, s5_91_fas, s5_92_facout, s5_92_fas, s5_100_facout, s5_100_fas, s5_101_facout, s5_101_fas, s5_102_facout, s5_102_fas, s5_110_facout, s5_110_fas, s5_111_facout, s5_111_fas, s5_112_facout, s5_112_fas, s5_120_facout, s5_120_fas, s5_121_facout, s5_121_fas, s5_122_facout, s5_122_fas, s5_130_facout, s5_130_fas, s5_131_facout, s5_131_fas, s5_132_facout, s5_132_fas, s5_140_facout, s5_140_fas, s5_141_facout, s5_141_fas, s5_142_facout, s5_142_fas, s5_150_facout, s5_150_fas, s5_151_facout, s5_151_fas, s5_152_facout, s5_152_fas, s5_160_facout, s5_160_fas, s5_161_facout, s5_161_fas, s5_162_facout, s5_162_fas, s5_170_facout, s5_170_fas, s5_171_facout, s5_171_fas, s5_172_facout, s5_172_fas, s5_180_facout, s5_180_fas, s5_181_facout, s5_181_fas, s5_182_facout, s5_182_fas, s5_190_facout, s5_190_fas, s5_191_facout, s5_191_fas, s5_192_facout, s5_192_fas, s5_200_facout, s5_200_fas, s5_201_facout, s5_201_fas, s5_202_facout, s5_202_fas, s5_210_facout, s5_210_fas, s5_211_facout, s5_211_fas, s5_212_facout, s5_212_fas, s5_220_facout, s5_220_fas, s5_221_facout, s5_221_fas, s5_222_facout, s5_222_fas, s5_230_facout, s5_230_fas, s5_231_facout, s5_231_fas, s5_232_facout, s5_232_fas, s5_240_facout, s5_240_fas, s5_241_facout, s5_241_fas, s5_242_facout, s5_242_fas, s5_250_facout, s5_250_fas, s5_251_facout, s5_251_fas, s5_252_facout, s5_252_fas, s5_260_facout, s5_260_fas, s5_261_facout, s5_261_fas, s5_262_facout, s5_262_fas, s5_270_facout, s5_270_fas, s5_271_facout, s5_271_fas, s5_272_facout, s5_272_fas, s5_280_facout, s5_280_fas, s5_281_facout, s5_281_fas, s5_282_facout, s5_282_fas, s5_290_facout, s5_290_fas, s5_291_facout, s5_291_fas, s5_292_facout, s5_292_fas, s5_300_facout, s5_300_fas, s5_301_facout, s5_301_fas, s5_302_facout, s5_302_fas, s5_310_facout, s5_310_fas, s5_311_facout, s5_311_fas, s5_312_facout, s5_312_fas, s5_320_facout, s5_320_fas, s5_321_facout, s5_321_fas, s5_322_facout, s5_322_fas, s5_330_facout, s5_330_fas, s5_331_facout, s5_331_fas, s5_332_facout, s5_332_fas, s5_340_facout, s5_340_fas, s5_341_facout, s5_341_fas, s5_342_facout, s5_342_fas, s5_350_facout, s5_350_fas, s5_351_facout, s5_351_fas, s5_352_facout, s5_352_fas, s5_360_facout, s5_360_fas, s5_361_facout, s5_361_fas, s5_362_facout, s5_362_fas, s5_370_facout, s5_370_fas, s5_371_facout, s5_371_fas, s5_372_facout, s5_372_fas, s5_380_facout, s5_380_fas, s5_381_facout, s5_381_fas, s5_382_facout, s5_382_fas, s5_390_facout, s5_390_fas, s5_391_facout, s5_391_fas, s5_392_facout, s5_392_fas, s5_400_facout, s5_400_fas, s5_401_facout, s5_401_fas, s5_402_facout, s5_402_fas, s5_410_facout, s5_410_fas, s5_411_facout, s5_411_fas, s5_412_facout, s5_412_fas, s5_420_facout, s5_420_fas, s5_421_facout, s5_421_fas, s5_422_facout, s5_422_fas, s5_430_facout, s5_430_fas, s5_431_facout, s5_431_fas, s5_432_facout, s5_432_fas, s5_440_facout, s5_440_fas, s5_441_facout, s5_441_fas, s5_442_facout, s5_442_fas, s5_450_facout, s5_450_fas, s5_451_facout, s5_451_fas, s5_452_facout, s5_452_fas, s5_460_facout, s5_460_fas, s5_461_facout, s5_461_fas, s5_462_facout, s5_462_fas, s5_470_facout, s5_470_fas, s5_471_facout, s5_471_fas, s5_472_facout, s5_472_fas, s5_480_facout, s5_480_fas, s5_481_facout, s5_481_fas, s5_482_facout, s5_482_fas, s5_490_facout, s5_490_fas, s5_491_facout, s5_491_fas, s5_492_facout, s5_492_fas, s5_500_facout, s5_500_fas, s5_501_facout, s5_501_fas, s5_502_facout, s5_502_fas, s5_510_facout, s5_510_fas, s5_511_facout, s5_511_fas, s5_512_facout, s5_512_fas, s5_520_facout, s5_520_fas, s5_521_facout, s5_521_fas, s5_522_facout, s5_522_fas, s5_530_facout, s5_530_fas, s5_531_facout, s5_531_fas, s5_532_facout, s5_532_fas, s5_540_facout, s5_540_fas, s5_541_facout, s5_541_fas, s5_542_facout, s5_542_fas, s5_550_facout, s5_550_fas, s5_551_facout, s5_551_fas, s5_552_facout, s5_552_fas, s5_560_facout, s5_560_fas, s5_561_facout, s5_561_fas, s5_570_facout, s5_570_fas;
/* ========================= Stage 5 ========================= */
half_adder s5_6ha0 ( .A(ps_66), .B(ps_65), .S(s5_60_has), .Cout(s5_60_hacout));
full_adder s5_7fa0 ( .A(ps_77), .B(ps_76), .Cin(ps_75), .S(s5_70_fas), .Cout(s5_70_facout));
half_adder s5_7ha0 ( .A(ps_74), .B(ps_73), .S(s5_70_has), .Cout(s5_70_hacout));
full_adder s5_8fa0 ( .A(ps_88), .B(ps_87), .Cin(ps_86), .S(s5_80_fas), .Cout(s5_80_facout));
full_adder s5_8fa1 ( .A(ps_85), .B(ps_84), .Cin(ps_83), .S(s5_81_fas), .Cout(s5_81_facout));
half_adder s5_8ha0 ( .A(ps_82), .B(ps_81), .S(s5_80_has), .Cout(s5_80_hacout));
full_adder s5_9fa0 ( .A(ps_97), .B(ps_96), .Cin(ps_95), .S(s5_90_fas), .Cout(s5_90_facout));
full_adder s5_9fa1 ( .A(ps_94), .B(ps_93), .Cin(ps_92), .S(s5_91_fas), .Cout(s5_91_facout));
full_adder s5_9fa2 ( .A(ps_91), .B(ps_90), .Cin(s4_90_has), .S(s5_92_fas), .Cout(s5_92_facout));
full_adder s5_10fa0 ( .A(ps_105), .B(ps_104), .Cin(ps_103), .S(s5_100_fas), .Cout(s5_100_facout));
full_adder s5_10fa1 ( .A(ps_102), .B(ps_101), .Cin(ps_100), .S(s5_101_fas), .Cout(s5_101_facout));
full_adder s5_10fa2 ( .A(s4_90_hacout), .B(s4_100_fas), .Cin(s4_100_has), .S(s5_102_fas), .Cout(s5_102_facout));
full_adder s5_11fa0 ( .A(ps_113), .B(ps_112), .Cin(ps_111), .S(s5_110_fas), .Cout(s5_110_facout));
full_adder s5_11fa1 ( .A(ps_110), .B(s4_100_facout), .Cin(s4_100_hacout), .S(s5_111_fas), .Cout(s5_111_facout));
full_adder s5_11fa2 ( .A(s4_110_fas), .B(s4_111_fas), .Cin(s4_110_has), .S(s5_112_fas), .Cout(s5_112_facout));
full_adder s5_12fa0 ( .A(ps_121), .B(ps_120), .Cin(s4_110_facout), .S(s5_120_fas), .Cout(s5_120_facout));
full_adder s5_12fa1 ( .A(s4_111_facout), .B(s4_110_hacout), .Cin(s4_120_fas), .S(s5_121_fas), .Cout(s5_121_facout));
full_adder s5_12fa2 ( .A(s4_121_fas), .B(s4_122_fas), .Cin(s4_120_has), .S(s5_122_fas), .Cout(s5_122_facout));
full_adder s5_13fa0 ( .A(s3_130_has), .B(s4_120_facout), .Cin(s4_121_facout), .S(s5_130_fas), .Cout(s5_130_facout));
full_adder s5_13fa1 ( .A(s4_122_facout), .B(s4_120_hacout), .Cin(s4_130_fas), .S(s5_131_fas), .Cout(s5_131_facout));
full_adder s5_13fa2 ( .A(s4_131_fas), .B(s4_132_fas), .Cin(s4_133_fas), .S(s5_132_fas), .Cout(s5_132_facout));
full_adder s5_14fa0 ( .A(s3_140_has), .B(s4_130_facout), .Cin(s4_131_facout), .S(s5_140_fas), .Cout(s5_140_facout));
full_adder s5_14fa1 ( .A(s4_132_facout), .B(s4_133_facout), .Cin(s4_140_fas), .S(s5_141_fas), .Cout(s5_141_facout));
full_adder s5_14fa2 ( .A(s4_141_fas), .B(s4_142_fas), .Cin(s4_143_fas), .S(s5_142_fas), .Cout(s5_142_facout));
full_adder s5_15fa0 ( .A(s3_150_has), .B(s4_140_facout), .Cin(s4_141_facout), .S(s5_150_fas), .Cout(s5_150_facout));
full_adder s5_15fa1 ( .A(s4_142_facout), .B(s4_143_facout), .Cin(s4_150_fas), .S(s5_151_fas), .Cout(s5_151_facout));
full_adder s5_15fa2 ( .A(s4_151_fas), .B(s4_152_fas), .Cin(s4_153_fas), .S(s5_152_fas), .Cout(s5_152_facout));
full_adder s5_16fa0 ( .A(s3_160_has), .B(s4_150_facout), .Cin(s4_151_facout), .S(s5_160_fas), .Cout(s5_160_facout));
full_adder s5_16fa1 ( .A(s4_152_facout), .B(s4_153_facout), .Cin(s4_160_fas), .S(s5_161_fas), .Cout(s5_161_facout));
full_adder s5_16fa2 ( .A(s4_161_fas), .B(s4_162_fas), .Cin(s4_163_fas), .S(s5_162_fas), .Cout(s5_162_facout));
full_adder s5_17fa0 ( .A(s3_170_has), .B(s4_160_facout), .Cin(s4_161_facout), .S(s5_170_fas), .Cout(s5_170_facout));
full_adder s5_17fa1 ( .A(s4_162_facout), .B(s4_163_facout), .Cin(s4_170_fas), .S(s5_171_fas), .Cout(s5_171_facout));
full_adder s5_17fa2 ( .A(s4_171_fas), .B(s4_172_fas), .Cin(s4_173_fas), .S(s5_172_fas), .Cout(s5_172_facout));
full_adder s5_18fa0 ( .A(s3_180_has), .B(s4_170_facout), .Cin(s4_171_facout), .S(s5_180_fas), .Cout(s5_180_facout));
full_adder s5_18fa1 ( .A(s4_172_facout), .B(s4_173_facout), .Cin(s4_180_fas), .S(s5_181_fas), .Cout(s5_181_facout));
full_adder s5_18fa2 ( .A(s4_181_fas), .B(s4_182_fas), .Cin(s4_183_fas), .S(s5_182_fas), .Cout(s5_182_facout));
full_adder s5_19fa0 ( .A(s3_195_fas), .B(s4_180_facout), .Cin(s4_181_facout), .S(s5_190_fas), .Cout(s5_190_facout));
full_adder s5_19fa1 ( .A(s4_182_facout), .B(s4_183_facout), .Cin(s4_190_fas), .S(s5_191_fas), .Cout(s5_191_facout));
full_adder s5_19fa2 ( .A(s4_191_fas), .B(s4_192_fas), .Cin(s4_193_fas), .S(s5_192_fas), .Cout(s5_192_facout));
full_adder s5_20fa0 ( .A(s3_205_fas), .B(s4_190_facout), .Cin(s4_191_facout), .S(s5_200_fas), .Cout(s5_200_facout));
full_adder s5_20fa1 ( .A(s4_192_facout), .B(s4_193_facout), .Cin(s4_200_fas), .S(s5_201_fas), .Cout(s5_201_facout));
full_adder s5_20fa2 ( .A(s4_201_fas), .B(s4_202_fas), .Cin(s4_203_fas), .S(s5_202_fas), .Cout(s5_202_facout));
full_adder s5_21fa0 ( .A(s3_215_fas), .B(s4_200_facout), .Cin(s4_201_facout), .S(s5_210_fas), .Cout(s5_210_facout));
full_adder s5_21fa1 ( .A(s4_202_facout), .B(s4_203_facout), .Cin(s4_210_fas), .S(s5_211_fas), .Cout(s5_211_facout));
full_adder s5_21fa2 ( .A(s4_211_fas), .B(s4_212_fas), .Cin(s4_213_fas), .S(s5_212_fas), .Cout(s5_212_facout));
full_adder s5_22fa0 ( .A(s3_225_fas), .B(s4_210_facout), .Cin(s4_211_facout), .S(s5_220_fas), .Cout(s5_220_facout));
full_adder s5_22fa1 ( .A(s4_212_facout), .B(s4_213_facout), .Cin(s4_220_fas), .S(s5_221_fas), .Cout(s5_221_facout));
full_adder s5_22fa2 ( .A(s4_221_fas), .B(s4_222_fas), .Cin(s4_223_fas), .S(s5_222_fas), .Cout(s5_222_facout));
full_adder s5_23fa0 ( .A(s3_235_fas), .B(s4_220_facout), .Cin(s4_221_facout), .S(s5_230_fas), .Cout(s5_230_facout));
full_adder s5_23fa1 ( .A(s4_222_facout), .B(s4_223_facout), .Cin(s4_230_fas), .S(s5_231_fas), .Cout(s5_231_facout));
full_adder s5_23fa2 ( .A(s4_231_fas), .B(s4_232_fas), .Cin(s4_233_fas), .S(s5_232_fas), .Cout(s5_232_facout));
full_adder s5_24fa0 ( .A(s3_245_fas), .B(s4_230_facout), .Cin(s4_231_facout), .S(s5_240_fas), .Cout(s5_240_facout));
full_adder s5_24fa1 ( .A(s4_232_facout), .B(s4_233_facout), .Cin(s4_240_fas), .S(s5_241_fas), .Cout(s5_241_facout));
full_adder s5_24fa2 ( .A(s4_241_fas), .B(s4_242_fas), .Cin(s4_243_fas), .S(s5_242_fas), .Cout(s5_242_facout));
full_adder s5_25fa0 ( .A(s3_255_fas), .B(s4_240_facout), .Cin(s4_241_facout), .S(s5_250_fas), .Cout(s5_250_facout));
full_adder s5_25fa1 ( .A(s4_242_facout), .B(s4_243_facout), .Cin(s4_250_fas), .S(s5_251_fas), .Cout(s5_251_facout));
full_adder s5_25fa2 ( .A(s4_251_fas), .B(s4_252_fas), .Cin(s4_253_fas), .S(s5_252_fas), .Cout(s5_252_facout));
full_adder s5_26fa0 ( .A(s3_265_fas), .B(s4_250_facout), .Cin(s4_251_facout), .S(s5_260_fas), .Cout(s5_260_facout));
full_adder s5_26fa1 ( .A(s4_252_facout), .B(s4_253_facout), .Cin(s4_260_fas), .S(s5_261_fas), .Cout(s5_261_facout));
full_adder s5_26fa2 ( .A(s4_261_fas), .B(s4_262_fas), .Cin(s4_263_fas), .S(s5_262_fas), .Cout(s5_262_facout));
full_adder s5_27fa0 ( .A(s3_275_fas), .B(s4_260_facout), .Cin(s4_261_facout), .S(s5_270_fas), .Cout(s5_270_facout));
full_adder s5_27fa1 ( .A(s4_262_facout), .B(s4_263_facout), .Cin(s4_270_fas), .S(s5_271_fas), .Cout(s5_271_facout));
full_adder s5_27fa2 ( .A(s4_271_fas), .B(s4_272_fas), .Cin(s4_273_fas), .S(s5_272_fas), .Cout(s5_272_facout));
full_adder s5_28fa0 ( .A(s3_285_fas), .B(s4_270_facout), .Cin(s4_271_facout), .S(s5_280_fas), .Cout(s5_280_facout));
full_adder s5_28fa1 ( .A(s4_272_facout), .B(s4_273_facout), .Cin(s4_280_fas), .S(s5_281_fas), .Cout(s5_281_facout));
full_adder s5_28fa2 ( .A(s4_281_fas), .B(s4_282_fas), .Cin(s4_283_fas), .S(s5_282_fas), .Cout(s5_282_facout));
full_adder s5_29fa0 ( .A(s3_295_fas), .B(s4_280_facout), .Cin(s4_281_facout), .S(s5_290_fas), .Cout(s5_290_facout));
full_adder s5_29fa1 ( .A(s4_282_facout), .B(s4_283_facout), .Cin(s4_290_fas), .S(s5_291_fas), .Cout(s5_291_facout));
full_adder s5_29fa2 ( .A(s4_291_fas), .B(s4_292_fas), .Cin(s4_293_fas), .S(s5_292_fas), .Cout(s5_292_facout));
full_adder s5_30fa0 ( .A(s3_305_fas), .B(s4_290_facout), .Cin(s4_291_facout), .S(s5_300_fas), .Cout(s5_300_facout));
full_adder s5_30fa1 ( .A(s4_292_facout), .B(s4_293_facout), .Cin(s4_300_fas), .S(s5_301_fas), .Cout(s5_301_facout));
full_adder s5_30fa2 ( .A(s4_301_fas), .B(s4_302_fas), .Cin(s4_303_fas), .S(s5_302_fas), .Cout(s5_302_facout));
full_adder s5_31fa0 ( .A(s3_315_fas), .B(s4_300_facout), .Cin(s4_301_facout), .S(s5_310_fas), .Cout(s5_310_facout));
full_adder s5_31fa1 ( .A(s4_302_facout), .B(s4_303_facout), .Cin(s4_310_fas), .S(s5_311_fas), .Cout(s5_311_facout));
full_adder s5_31fa2 ( .A(s4_311_fas), .B(s4_312_fas), .Cin(s4_313_fas), .S(s5_312_fas), .Cout(s5_312_facout));
full_adder s5_32fa0 ( .A(s3_325_fas), .B(s4_310_facout), .Cin(s4_311_facout), .S(s5_320_fas), .Cout(s5_320_facout));
full_adder s5_32fa1 ( .A(s4_312_facout), .B(s4_313_facout), .Cin(s4_320_fas), .S(s5_321_fas), .Cout(s5_321_facout));
full_adder s5_32fa2 ( .A(s4_321_fas), .B(s4_322_fas), .Cin(s4_323_fas), .S(s5_322_fas), .Cout(s5_322_facout));
full_adder s5_33fa0 ( .A(s3_335_fas), .B(s4_320_facout), .Cin(s4_321_facout), .S(s5_330_fas), .Cout(s5_330_facout));
full_adder s5_33fa1 ( .A(s4_322_facout), .B(s4_323_facout), .Cin(s4_330_fas), .S(s5_331_fas), .Cout(s5_331_facout));
full_adder s5_33fa2 ( .A(s4_331_fas), .B(s4_332_fas), .Cin(s4_333_fas), .S(s5_332_fas), .Cout(s5_332_facout));
full_adder s5_34fa0 ( .A(s3_345_fas), .B(s4_330_facout), .Cin(s4_331_facout), .S(s5_340_fas), .Cout(s5_340_facout));
full_adder s5_34fa1 ( .A(s4_332_facout), .B(s4_333_facout), .Cin(s4_340_fas), .S(s5_341_fas), .Cout(s5_341_facout));
full_adder s5_34fa2 ( .A(s4_341_fas), .B(s4_342_fas), .Cin(s4_343_fas), .S(s5_342_fas), .Cout(s5_342_facout));
full_adder s5_35fa0 ( .A(s3_355_fas), .B(s4_340_facout), .Cin(s4_341_facout), .S(s5_350_fas), .Cout(s5_350_facout));
full_adder s5_35fa1 ( .A(s4_342_facout), .B(s4_343_facout), .Cin(s4_350_fas), .S(s5_351_fas), .Cout(s5_351_facout));
full_adder s5_35fa2 ( .A(s4_351_fas), .B(s4_352_fas), .Cin(s4_353_fas), .S(s5_352_fas), .Cout(s5_352_facout));
full_adder s5_36fa0 ( .A(s3_365_fas), .B(s4_350_facout), .Cin(s4_351_facout), .S(s5_360_fas), .Cout(s5_360_facout));
full_adder s5_36fa1 ( .A(s4_352_facout), .B(s4_353_facout), .Cin(s4_360_fas), .S(s5_361_fas), .Cout(s5_361_facout));
full_adder s5_36fa2 ( .A(s4_361_fas), .B(s4_362_fas), .Cin(s4_363_fas), .S(s5_362_fas), .Cout(s5_362_facout));
full_adder s5_37fa0 ( .A(s3_375_fas), .B(s4_360_facout), .Cin(s4_361_facout), .S(s5_370_fas), .Cout(s5_370_facout));
full_adder s5_37fa1 ( .A(s4_362_facout), .B(s4_363_facout), .Cin(s4_370_fas), .S(s5_371_fas), .Cout(s5_371_facout));
full_adder s5_37fa2 ( .A(s4_371_fas), .B(s4_372_fas), .Cin(s4_373_fas), .S(s5_372_fas), .Cout(s5_372_facout));
full_adder s5_38fa0 ( .A(s3_385_fas), .B(s4_370_facout), .Cin(s4_371_facout), .S(s5_380_fas), .Cout(s5_380_facout));
full_adder s5_38fa1 ( .A(s4_372_facout), .B(s4_373_facout), .Cin(s4_380_fas), .S(s5_381_fas), .Cout(s5_381_facout));
full_adder s5_38fa2 ( .A(s4_381_fas), .B(s4_382_fas), .Cin(s4_383_fas), .S(s5_382_fas), .Cout(s5_382_facout));
full_adder s5_39fa0 ( .A(s3_395_fas), .B(s4_380_facout), .Cin(s4_381_facout), .S(s5_390_fas), .Cout(s5_390_facout));
full_adder s5_39fa1 ( .A(s4_382_facout), .B(s4_383_facout), .Cin(s4_390_fas), .S(s5_391_fas), .Cout(s5_391_facout));
full_adder s5_39fa2 ( .A(s4_391_fas), .B(s4_392_fas), .Cin(s4_393_fas), .S(s5_392_fas), .Cout(s5_392_facout));
full_adder s5_40fa0 ( .A(s3_405_fas), .B(s4_390_facout), .Cin(s4_391_facout), .S(s5_400_fas), .Cout(s5_400_facout));
full_adder s5_40fa1 ( .A(s4_392_facout), .B(s4_393_facout), .Cin(s4_400_fas), .S(s5_401_fas), .Cout(s5_401_facout));
full_adder s5_40fa2 ( .A(s4_401_fas), .B(s4_402_fas), .Cin(s4_403_fas), .S(s5_402_fas), .Cout(s5_402_facout));
full_adder s5_41fa0 ( .A(s3_415_fas), .B(s4_400_facout), .Cin(s4_401_facout), .S(s5_410_fas), .Cout(s5_410_facout));
full_adder s5_41fa1 ( .A(s4_402_facout), .B(s4_403_facout), .Cin(s4_410_fas), .S(s5_411_fas), .Cout(s5_411_facout));
full_adder s5_41fa2 ( .A(s4_411_fas), .B(s4_412_fas), .Cin(s4_413_fas), .S(s5_412_fas), .Cout(s5_412_facout));
full_adder s5_42fa0 ( .A(s3_425_fas), .B(s4_410_facout), .Cin(s4_411_facout), .S(s5_420_fas), .Cout(s5_420_facout));
full_adder s5_42fa1 ( .A(s4_412_facout), .B(s4_413_facout), .Cin(s4_420_fas), .S(s5_421_fas), .Cout(s5_421_facout));
full_adder s5_42fa2 ( .A(s4_421_fas), .B(s4_422_fas), .Cin(s4_423_fas), .S(s5_422_fas), .Cout(s5_422_facout));
full_adder s5_43fa0 ( .A(s3_435_fas), .B(s4_420_facout), .Cin(s4_421_facout), .S(s5_430_fas), .Cout(s5_430_facout));
full_adder s5_43fa1 ( .A(s4_422_facout), .B(s4_423_facout), .Cin(s4_430_fas), .S(s5_431_fas), .Cout(s5_431_facout));
full_adder s5_43fa2 ( .A(s4_431_fas), .B(s4_432_fas), .Cin(s4_433_fas), .S(s5_432_fas), .Cout(s5_432_facout));
full_adder s5_44fa0 ( .A(s3_445_fas), .B(s4_430_facout), .Cin(s4_431_facout), .S(s5_440_fas), .Cout(s5_440_facout));
full_adder s5_44fa1 ( .A(s4_432_facout), .B(s4_433_facout), .Cin(s4_440_fas), .S(s5_441_fas), .Cout(s5_441_facout));
full_adder s5_44fa2 ( .A(s4_441_fas), .B(s4_442_fas), .Cin(s4_443_fas), .S(s5_442_fas), .Cout(s5_442_facout));
full_adder s5_45fa0 ( .A(s3_455_fas), .B(s4_440_facout), .Cin(s4_441_facout), .S(s5_450_fas), .Cout(s5_450_facout));
full_adder s5_45fa1 ( .A(s4_442_facout), .B(s4_443_facout), .Cin(s4_450_fas), .S(s5_451_fas), .Cout(s5_451_facout));
full_adder s5_45fa2 ( .A(s4_451_fas), .B(s4_452_fas), .Cin(s4_453_fas), .S(s5_452_fas), .Cout(s5_452_facout));
full_adder s5_46fa0 ( .A(s3_464_fas), .B(s4_450_facout), .Cin(s4_451_facout), .S(s5_460_fas), .Cout(s5_460_facout));
full_adder s5_46fa1 ( .A(s4_452_facout), .B(s4_453_facout), .Cin(s4_460_fas), .S(s5_461_fas), .Cout(s5_461_facout));
full_adder s5_46fa2 ( .A(s4_461_fas), .B(s4_462_fas), .Cin(s4_463_fas), .S(s5_462_fas), .Cout(s5_462_facout));
full_adder s5_47fa0 ( .A(s3_473_fas), .B(s4_460_facout), .Cin(s4_461_facout), .S(s5_470_fas), .Cout(s5_470_facout));
full_adder s5_47fa1 ( .A(s4_462_facout), .B(s4_463_facout), .Cin(s4_470_fas), .S(s5_471_fas), .Cout(s5_471_facout));
full_adder s5_47fa2 ( .A(s4_471_fas), .B(s4_472_fas), .Cin(s4_473_fas), .S(s5_472_fas), .Cout(s5_472_facout));
full_adder s5_48fa0 ( .A(s3_482_fas), .B(s4_470_facout), .Cin(s4_471_facout), .S(s5_480_fas), .Cout(s5_480_facout));
full_adder s5_48fa1 ( .A(s4_472_facout), .B(s4_473_facout), .Cin(s4_480_fas), .S(s5_481_fas), .Cout(s5_481_facout));
full_adder s5_48fa2 ( .A(s4_481_fas), .B(s4_482_fas), .Cin(s4_483_fas), .S(s5_482_fas), .Cout(s5_482_facout));
full_adder s5_49fa0 ( .A(s3_491_fas), .B(s4_480_facout), .Cin(s4_481_facout), .S(s5_490_fas), .Cout(s5_490_facout));
full_adder s5_49fa1 ( .A(s4_482_facout), .B(s4_483_facout), .Cin(s4_490_fas), .S(s5_491_fas), .Cout(s5_491_facout));
full_adder s5_49fa2 ( .A(s4_491_fas), .B(s4_492_fas), .Cin(s4_493_fas), .S(s5_492_fas), .Cout(s5_492_facout));
full_adder s5_50fa0 ( .A(s3_500_fas), .B(s4_490_facout), .Cin(s4_491_facout), .S(s5_500_fas), .Cout(s5_500_facout));
full_adder s5_50fa1 ( .A(s4_492_facout), .B(s4_493_facout), .Cin(s4_500_fas), .S(s5_501_fas), .Cout(s5_501_facout));
full_adder s5_50fa2 ( .A(s4_501_fas), .B(s4_502_fas), .Cin(s4_503_fas), .S(s5_502_fas), .Cout(s5_502_facout));
full_adder s5_51fa0 ( .A(s3_500_facout), .B(s4_500_facout), .Cin(s4_501_facout), .S(s5_510_fas), .Cout(s5_510_facout));
full_adder s5_51fa1 ( .A(s4_502_facout), .B(s4_503_facout), .Cin(s4_510_fas), .S(s5_511_fas), .Cout(s5_511_facout));
full_adder s5_51fa2 ( .A(s4_511_fas), .B(s4_512_fas), .Cin(s4_513_fas), .S(s5_512_fas), .Cout(s5_512_facout));
full_adder s5_52fa0 ( .A(ps_5222), .B(ps_5221), .Cin(s4_510_facout), .S(s5_520_fas), .Cout(s5_520_facout));
full_adder s5_52fa1 ( .A(s4_511_facout), .B(s4_512_facout), .Cin(s4_513_facout), .S(s5_521_fas), .Cout(s5_521_facout));
full_adder s5_52fa2 ( .A(s4_520_fas), .B(s4_521_fas), .Cin(s4_522_fas), .S(s5_522_fas), .Cout(s5_522_facout));
full_adder s5_53fa0 ( .A(ps_5325), .B(ps_5324), .Cin(ps_5323), .S(s5_530_fas), .Cout(s5_530_facout));
full_adder s5_53fa1 ( .A(ps_5322), .B(s4_520_facout), .Cin(s4_521_facout), .S(s5_531_fas), .Cout(s5_531_facout));
full_adder s5_53fa2 ( .A(s4_522_facout), .B(s4_530_fas), .Cin(s4_531_fas), .S(s5_532_fas), .Cout(s5_532_facout));
full_adder s5_54fa0 ( .A(ps_5428), .B(ps_5427), .Cin(ps_5426), .S(s5_540_fas), .Cout(s5_540_facout));
full_adder s5_54fa1 ( .A(ps_5425), .B(ps_5424), .Cin(ps_5423), .S(s5_541_fas), .Cout(s5_541_facout));
full_adder s5_54fa2 ( .A(s4_530_facout), .B(s4_531_facout), .Cin(s4_540_fas), .S(s5_542_fas), .Cout(s5_542_facout));
full_adder s5_55fa0 ( .A(ps_5531), .B(ps_5530), .Cin(ps_5529), .S(s5_550_fas), .Cout(s5_550_facout));
full_adder s5_55fa1 ( .A(ps_5528), .B(ps_5527), .Cin(ps_5526), .S(s5_551_fas), .Cout(s5_551_facout));
full_adder s5_55fa2 ( .A(ps_5525), .B(ps_5524), .Cin(s4_540_facout), .S(s5_552_fas), .Cout(s5_552_facout));
full_adder s5_56fa0 ( .A(ps_5631), .B(ps_5630), .Cin(ps_5629), .S(s5_560_fas), .Cout(s5_560_facout));
full_adder s5_56fa1 ( .A(ps_5628), .B(ps_5627), .Cin(ps_5626), .S(s5_561_fas), .Cout(s5_561_facout));
full_adder s5_57fa0 ( .A(ps_5731), .B(ps_5730), .Cin(ps_5729), .S(s5_570_fas), .Cout(s5_570_facout));
logic s6_40_hacout, s6_40_has, s6_50_facout, s6_50_fas, s6_50_hacout, s6_50_has, s6_60_facout, s6_60_fas, s6_61_facout, s6_61_fas, s6_70_facout, s6_70_fas, s6_71_facout, s6_71_fas, s6_80_facout, s6_80_fas, s6_81_facout, s6_81_fas, s6_90_facout, s6_90_fas, s6_91_facout, s6_91_fas, s6_100_facout, s6_100_fas, s6_101_facout, s6_101_fas, s6_110_facout, s6_110_fas, s6_111_facout, s6_111_fas, s6_120_facout, s6_120_fas, s6_121_facout, s6_121_fas, s6_130_facout, s6_130_fas, s6_131_facout, s6_131_fas, s6_140_facout, s6_140_fas, s6_141_facout, s6_141_fas, s6_150_facout, s6_150_fas, s6_151_facout, s6_151_fas, s6_160_facout, s6_160_fas, s6_161_facout, s6_161_fas, s6_170_facout, s6_170_fas, s6_171_facout, s6_171_fas, s6_180_facout, s6_180_fas, s6_181_facout, s6_181_fas, s6_190_facout, s6_190_fas, s6_191_facout, s6_191_fas, s6_200_facout, s6_200_fas, s6_201_facout, s6_201_fas, s6_210_facout, s6_210_fas, s6_211_facout, s6_211_fas, s6_220_facout, s6_220_fas, s6_221_facout, s6_221_fas, s6_230_facout, s6_230_fas, s6_231_facout, s6_231_fas, s6_240_facout, s6_240_fas, s6_241_facout, s6_241_fas, s6_250_facout, s6_250_fas, s6_251_facout, s6_251_fas, s6_260_facout, s6_260_fas, s6_261_facout, s6_261_fas, s6_270_facout, s6_270_fas, s6_271_facout, s6_271_fas, s6_280_facout, s6_280_fas, s6_281_facout, s6_281_fas, s6_290_facout, s6_290_fas, s6_291_facout, s6_291_fas, s6_300_facout, s6_300_fas, s6_301_facout, s6_301_fas, s6_310_facout, s6_310_fas, s6_311_facout, s6_311_fas, s6_320_facout, s6_320_fas, s6_321_facout, s6_321_fas, s6_330_facout, s6_330_fas, s6_331_facout, s6_331_fas, s6_340_facout, s6_340_fas, s6_341_facout, s6_341_fas, s6_350_facout, s6_350_fas, s6_351_facout, s6_351_fas, s6_360_facout, s6_360_fas, s6_361_facout, s6_361_fas, s6_370_facout, s6_370_fas, s6_371_facout, s6_371_fas, s6_380_facout, s6_380_fas, s6_381_facout, s6_381_fas, s6_390_facout, s6_390_fas, s6_391_facout, s6_391_fas, s6_400_facout, s6_400_fas, s6_401_facout, s6_401_fas, s6_410_facout, s6_410_fas, s6_411_facout, s6_411_fas, s6_420_facout, s6_420_fas, s6_421_facout, s6_421_fas, s6_430_facout, s6_430_fas, s6_431_facout, s6_431_fas, s6_440_facout, s6_440_fas, s6_441_facout, s6_441_fas, s6_450_facout, s6_450_fas, s6_451_facout, s6_451_fas, s6_460_facout, s6_460_fas, s6_461_facout, s6_461_fas, s6_470_facout, s6_470_fas, s6_471_facout, s6_471_fas, s6_480_facout, s6_480_fas, s6_481_facout, s6_481_fas, s6_490_facout, s6_490_fas, s6_491_facout, s6_491_fas, s6_500_facout, s6_500_fas, s6_501_facout, s6_501_fas, s6_510_facout, s6_510_fas, s6_511_facout, s6_511_fas, s6_520_facout, s6_520_fas, s6_521_facout, s6_521_fas, s6_530_facout, s6_530_fas, s6_531_facout, s6_531_fas, s6_540_facout, s6_540_fas, s6_541_facout, s6_541_fas, s6_550_facout, s6_550_fas, s6_551_facout, s6_551_fas, s6_560_facout, s6_560_fas, s6_561_facout, s6_561_fas, s6_570_facout, s6_570_fas, s6_571_facout, s6_571_fas, s6_580_facout, s6_580_fas, s6_581_facout, s6_581_fas, s6_590_facout, s6_590_fas;
/* ========================= Stage 6 ========================= */
half_adder s6_4ha0 ( .A(ps_44), .B(ps_43), .S(s6_40_has), .Cout(s6_40_hacout));
full_adder s6_5fa0 ( .A(ps_55), .B(ps_54), .Cin(ps_53), .S(s6_50_fas), .Cout(s6_50_facout));
half_adder s6_5ha0 ( .A(ps_52), .B(ps_51), .S(s6_50_has), .Cout(s6_50_hacout));
full_adder s6_6fa0 ( .A(ps_64), .B(ps_63), .Cin(ps_62), .S(s6_60_fas), .Cout(s6_60_facout));
full_adder s6_6fa1 ( .A(ps_61), .B(ps_60), .Cin(s5_60_has), .S(s6_61_fas), .Cout(s6_61_facout));
full_adder s6_7fa0 ( .A(ps_72), .B(ps_71), .Cin(ps_70), .S(s6_70_fas), .Cout(s6_70_facout));
full_adder s6_7fa1 ( .A(s5_60_hacout), .B(s5_70_fas), .Cin(s5_70_has), .S(s6_71_fas), .Cout(s6_71_facout));
full_adder s6_8fa0 ( .A(ps_80), .B(s5_70_facout), .Cin(s5_70_hacout), .S(s6_80_fas), .Cout(s6_80_facout));
full_adder s6_8fa1 ( .A(s5_80_fas), .B(s5_81_fas), .Cin(s5_80_has), .S(s6_81_fas), .Cout(s6_81_facout));
full_adder s6_9fa0 ( .A(s5_80_facout), .B(s5_81_facout), .Cin(s5_80_hacout), .S(s6_90_fas), .Cout(s6_90_facout));
full_adder s6_9fa1 ( .A(s5_90_fas), .B(s5_91_fas), .Cin(s5_92_fas), .S(s6_91_fas), .Cout(s6_91_facout));
full_adder s6_10fa0 ( .A(s5_90_facout), .B(s5_91_facout), .Cin(s5_92_facout), .S(s6_100_fas), .Cout(s6_100_facout));
full_adder s6_10fa1 ( .A(s5_100_fas), .B(s5_101_fas), .Cin(s5_102_fas), .S(s6_101_fas), .Cout(s6_101_facout));
full_adder s6_11fa0 ( .A(s5_100_facout), .B(s5_101_facout), .Cin(s5_102_facout), .S(s6_110_fas), .Cout(s6_110_facout));
full_adder s6_11fa1 ( .A(s5_110_fas), .B(s5_111_fas), .Cin(s5_112_fas), .S(s6_111_fas), .Cout(s6_111_facout));
full_adder s6_12fa0 ( .A(s5_110_facout), .B(s5_111_facout), .Cin(s5_112_facout), .S(s6_120_fas), .Cout(s6_120_facout));
full_adder s6_12fa1 ( .A(s5_120_fas), .B(s5_121_fas), .Cin(s5_122_fas), .S(s6_121_fas), .Cout(s6_121_facout));
full_adder s6_13fa0 ( .A(s5_120_facout), .B(s5_121_facout), .Cin(s5_122_facout), .S(s6_130_fas), .Cout(s6_130_facout));
full_adder s6_13fa1 ( .A(s5_130_fas), .B(s5_131_fas), .Cin(s5_132_fas), .S(s6_131_fas), .Cout(s6_131_facout));
full_adder s6_14fa0 ( .A(s5_130_facout), .B(s5_131_facout), .Cin(s5_132_facout), .S(s6_140_fas), .Cout(s6_140_facout));
full_adder s6_14fa1 ( .A(s5_140_fas), .B(s5_141_fas), .Cin(s5_142_fas), .S(s6_141_fas), .Cout(s6_141_facout));
full_adder s6_15fa0 ( .A(s5_140_facout), .B(s5_141_facout), .Cin(s5_142_facout), .S(s6_150_fas), .Cout(s6_150_facout));
full_adder s6_15fa1 ( .A(s5_150_fas), .B(s5_151_fas), .Cin(s5_152_fas), .S(s6_151_fas), .Cout(s6_151_facout));
full_adder s6_16fa0 ( .A(s5_150_facout), .B(s5_151_facout), .Cin(s5_152_facout), .S(s6_160_fas), .Cout(s6_160_facout));
full_adder s6_16fa1 ( .A(s5_160_fas), .B(s5_161_fas), .Cin(s5_162_fas), .S(s6_161_fas), .Cout(s6_161_facout));
full_adder s6_17fa0 ( .A(s5_160_facout), .B(s5_161_facout), .Cin(s5_162_facout), .S(s6_170_fas), .Cout(s6_170_facout));
full_adder s6_17fa1 ( .A(s5_170_fas), .B(s5_171_fas), .Cin(s5_172_fas), .S(s6_171_fas), .Cout(s6_171_facout));
full_adder s6_18fa0 ( .A(s5_170_facout), .B(s5_171_facout), .Cin(s5_172_facout), .S(s6_180_fas), .Cout(s6_180_facout));
full_adder s6_18fa1 ( .A(s5_180_fas), .B(s5_181_fas), .Cin(s5_182_fas), .S(s6_181_fas), .Cout(s6_181_facout));
full_adder s6_19fa0 ( .A(s5_180_facout), .B(s5_181_facout), .Cin(s5_182_facout), .S(s6_190_fas), .Cout(s6_190_facout));
full_adder s6_19fa1 ( .A(s5_190_fas), .B(s5_191_fas), .Cin(s5_192_fas), .S(s6_191_fas), .Cout(s6_191_facout));
full_adder s6_20fa0 ( .A(s5_190_facout), .B(s5_191_facout), .Cin(s5_192_facout), .S(s6_200_fas), .Cout(s6_200_facout));
full_adder s6_20fa1 ( .A(s5_200_fas), .B(s5_201_fas), .Cin(s5_202_fas), .S(s6_201_fas), .Cout(s6_201_facout));
full_adder s6_21fa0 ( .A(s5_200_facout), .B(s5_201_facout), .Cin(s5_202_facout), .S(s6_210_fas), .Cout(s6_210_facout));
full_adder s6_21fa1 ( .A(s5_210_fas), .B(s5_211_fas), .Cin(s5_212_fas), .S(s6_211_fas), .Cout(s6_211_facout));
full_adder s6_22fa0 ( .A(s5_210_facout), .B(s5_211_facout), .Cin(s5_212_facout), .S(s6_220_fas), .Cout(s6_220_facout));
full_adder s6_22fa1 ( .A(s5_220_fas), .B(s5_221_fas), .Cin(s5_222_fas), .S(s6_221_fas), .Cout(s6_221_facout));
full_adder s6_23fa0 ( .A(s5_220_facout), .B(s5_221_facout), .Cin(s5_222_facout), .S(s6_230_fas), .Cout(s6_230_facout));
full_adder s6_23fa1 ( .A(s5_230_fas), .B(s5_231_fas), .Cin(s5_232_fas), .S(s6_231_fas), .Cout(s6_231_facout));
full_adder s6_24fa0 ( .A(s5_230_facout), .B(s5_231_facout), .Cin(s5_232_facout), .S(s6_240_fas), .Cout(s6_240_facout));
full_adder s6_24fa1 ( .A(s5_240_fas), .B(s5_241_fas), .Cin(s5_242_fas), .S(s6_241_fas), .Cout(s6_241_facout));
full_adder s6_25fa0 ( .A(s5_240_facout), .B(s5_241_facout), .Cin(s5_242_facout), .S(s6_250_fas), .Cout(s6_250_facout));
full_adder s6_25fa1 ( .A(s5_250_fas), .B(s5_251_fas), .Cin(s5_252_fas), .S(s6_251_fas), .Cout(s6_251_facout));
full_adder s6_26fa0 ( .A(s5_250_facout), .B(s5_251_facout), .Cin(s5_252_facout), .S(s6_260_fas), .Cout(s6_260_facout));
full_adder s6_26fa1 ( .A(s5_260_fas), .B(s5_261_fas), .Cin(s5_262_fas), .S(s6_261_fas), .Cout(s6_261_facout));
full_adder s6_27fa0 ( .A(s5_260_facout), .B(s5_261_facout), .Cin(s5_262_facout), .S(s6_270_fas), .Cout(s6_270_facout));
full_adder s6_27fa1 ( .A(s5_270_fas), .B(s5_271_fas), .Cin(s5_272_fas), .S(s6_271_fas), .Cout(s6_271_facout));
full_adder s6_28fa0 ( .A(s5_270_facout), .B(s5_271_facout), .Cin(s5_272_facout), .S(s6_280_fas), .Cout(s6_280_facout));
full_adder s6_28fa1 ( .A(s5_280_fas), .B(s5_281_fas), .Cin(s5_282_fas), .S(s6_281_fas), .Cout(s6_281_facout));
full_adder s6_29fa0 ( .A(s5_280_facout), .B(s5_281_facout), .Cin(s5_282_facout), .S(s6_290_fas), .Cout(s6_290_facout));
full_adder s6_29fa1 ( .A(s5_290_fas), .B(s5_291_fas), .Cin(s5_292_fas), .S(s6_291_fas), .Cout(s6_291_facout));
full_adder s6_30fa0 ( .A(s5_290_facout), .B(s5_291_facout), .Cin(s5_292_facout), .S(s6_300_fas), .Cout(s6_300_facout));
full_adder s6_30fa1 ( .A(s5_300_fas), .B(s5_301_fas), .Cin(s5_302_fas), .S(s6_301_fas), .Cout(s6_301_facout));
full_adder s6_31fa0 ( .A(s5_300_facout), .B(s5_301_facout), .Cin(s5_302_facout), .S(s6_310_fas), .Cout(s6_310_facout));
full_adder s6_31fa1 ( .A(s5_310_fas), .B(s5_311_fas), .Cin(s5_312_fas), .S(s6_311_fas), .Cout(s6_311_facout));
full_adder s6_32fa0 ( .A(s5_310_facout), .B(s5_311_facout), .Cin(s5_312_facout), .S(s6_320_fas), .Cout(s6_320_facout));
full_adder s6_32fa1 ( .A(s5_320_fas), .B(s5_321_fas), .Cin(s5_322_fas), .S(s6_321_fas), .Cout(s6_321_facout));
full_adder s6_33fa0 ( .A(s5_320_facout), .B(s5_321_facout), .Cin(s5_322_facout), .S(s6_330_fas), .Cout(s6_330_facout));
full_adder s6_33fa1 ( .A(s5_330_fas), .B(s5_331_fas), .Cin(s5_332_fas), .S(s6_331_fas), .Cout(s6_331_facout));
full_adder s6_34fa0 ( .A(s5_330_facout), .B(s5_331_facout), .Cin(s5_332_facout), .S(s6_340_fas), .Cout(s6_340_facout));
full_adder s6_34fa1 ( .A(s5_340_fas), .B(s5_341_fas), .Cin(s5_342_fas), .S(s6_341_fas), .Cout(s6_341_facout));
full_adder s6_35fa0 ( .A(s5_340_facout), .B(s5_341_facout), .Cin(s5_342_facout), .S(s6_350_fas), .Cout(s6_350_facout));
full_adder s6_35fa1 ( .A(s5_350_fas), .B(s5_351_fas), .Cin(s5_352_fas), .S(s6_351_fas), .Cout(s6_351_facout));
full_adder s6_36fa0 ( .A(s5_350_facout), .B(s5_351_facout), .Cin(s5_352_facout), .S(s6_360_fas), .Cout(s6_360_facout));
full_adder s6_36fa1 ( .A(s5_360_fas), .B(s5_361_fas), .Cin(s5_362_fas), .S(s6_361_fas), .Cout(s6_361_facout));
full_adder s6_37fa0 ( .A(s5_360_facout), .B(s5_361_facout), .Cin(s5_362_facout), .S(s6_370_fas), .Cout(s6_370_facout));
full_adder s6_37fa1 ( .A(s5_370_fas), .B(s5_371_fas), .Cin(s5_372_fas), .S(s6_371_fas), .Cout(s6_371_facout));
full_adder s6_38fa0 ( .A(s5_370_facout), .B(s5_371_facout), .Cin(s5_372_facout), .S(s6_380_fas), .Cout(s6_380_facout));
full_adder s6_38fa1 ( .A(s5_380_fas), .B(s5_381_fas), .Cin(s5_382_fas), .S(s6_381_fas), .Cout(s6_381_facout));
full_adder s6_39fa0 ( .A(s5_380_facout), .B(s5_381_facout), .Cin(s5_382_facout), .S(s6_390_fas), .Cout(s6_390_facout));
full_adder s6_39fa1 ( .A(s5_390_fas), .B(s5_391_fas), .Cin(s5_392_fas), .S(s6_391_fas), .Cout(s6_391_facout));
full_adder s6_40fa0 ( .A(s5_390_facout), .B(s5_391_facout), .Cin(s5_392_facout), .S(s6_400_fas), .Cout(s6_400_facout));
full_adder s6_40fa1 ( .A(s5_400_fas), .B(s5_401_fas), .Cin(s5_402_fas), .S(s6_401_fas), .Cout(s6_401_facout));
full_adder s6_41fa0 ( .A(s5_400_facout), .B(s5_401_facout), .Cin(s5_402_facout), .S(s6_410_fas), .Cout(s6_410_facout));
full_adder s6_41fa1 ( .A(s5_410_fas), .B(s5_411_fas), .Cin(s5_412_fas), .S(s6_411_fas), .Cout(s6_411_facout));
full_adder s6_42fa0 ( .A(s5_410_facout), .B(s5_411_facout), .Cin(s5_412_facout), .S(s6_420_fas), .Cout(s6_420_facout));
full_adder s6_42fa1 ( .A(s5_420_fas), .B(s5_421_fas), .Cin(s5_422_fas), .S(s6_421_fas), .Cout(s6_421_facout));
full_adder s6_43fa0 ( .A(s5_420_facout), .B(s5_421_facout), .Cin(s5_422_facout), .S(s6_430_fas), .Cout(s6_430_facout));
full_adder s6_43fa1 ( .A(s5_430_fas), .B(s5_431_fas), .Cin(s5_432_fas), .S(s6_431_fas), .Cout(s6_431_facout));
full_adder s6_44fa0 ( .A(s5_430_facout), .B(s5_431_facout), .Cin(s5_432_facout), .S(s6_440_fas), .Cout(s6_440_facout));
full_adder s6_44fa1 ( .A(s5_440_fas), .B(s5_441_fas), .Cin(s5_442_fas), .S(s6_441_fas), .Cout(s6_441_facout));
full_adder s6_45fa0 ( .A(s5_440_facout), .B(s5_441_facout), .Cin(s5_442_facout), .S(s6_450_fas), .Cout(s6_450_facout));
full_adder s6_45fa1 ( .A(s5_450_fas), .B(s5_451_fas), .Cin(s5_452_fas), .S(s6_451_fas), .Cout(s6_451_facout));
full_adder s6_46fa0 ( .A(s5_450_facout), .B(s5_451_facout), .Cin(s5_452_facout), .S(s6_460_fas), .Cout(s6_460_facout));
full_adder s6_46fa1 ( .A(s5_460_fas), .B(s5_461_fas), .Cin(s5_462_fas), .S(s6_461_fas), .Cout(s6_461_facout));
full_adder s6_47fa0 ( .A(s5_460_facout), .B(s5_461_facout), .Cin(s5_462_facout), .S(s6_470_fas), .Cout(s6_470_facout));
full_adder s6_47fa1 ( .A(s5_470_fas), .B(s5_471_fas), .Cin(s5_472_fas), .S(s6_471_fas), .Cout(s6_471_facout));
full_adder s6_48fa0 ( .A(s5_470_facout), .B(s5_471_facout), .Cin(s5_472_facout), .S(s6_480_fas), .Cout(s6_480_facout));
full_adder s6_48fa1 ( .A(s5_480_fas), .B(s5_481_fas), .Cin(s5_482_fas), .S(s6_481_fas), .Cout(s6_481_facout));
full_adder s6_49fa0 ( .A(s5_480_facout), .B(s5_481_facout), .Cin(s5_482_facout), .S(s6_490_fas), .Cout(s6_490_facout));
full_adder s6_49fa1 ( .A(s5_490_fas), .B(s5_491_fas), .Cin(s5_492_fas), .S(s6_491_fas), .Cout(s6_491_facout));
full_adder s6_50fa0 ( .A(s5_490_facout), .B(s5_491_facout), .Cin(s5_492_facout), .S(s6_500_fas), .Cout(s6_500_facout));
full_adder s6_50fa1 ( .A(s5_500_fas), .B(s5_501_fas), .Cin(s5_502_fas), .S(s6_501_fas), .Cout(s6_501_facout));
full_adder s6_51fa0 ( .A(s5_500_facout), .B(s5_501_facout), .Cin(s5_502_facout), .S(s6_510_fas), .Cout(s6_510_facout));
full_adder s6_51fa1 ( .A(s5_510_fas), .B(s5_511_fas), .Cin(s5_512_fas), .S(s6_511_fas), .Cout(s6_511_facout));
full_adder s6_52fa0 ( .A(s5_510_facout), .B(s5_511_facout), .Cin(s5_512_facout), .S(s6_520_fas), .Cout(s6_520_facout));
full_adder s6_52fa1 ( .A(s5_520_fas), .B(s5_521_fas), .Cin(s5_522_fas), .S(s6_521_fas), .Cout(s6_521_facout));
full_adder s6_53fa0 ( .A(s5_520_facout), .B(s5_521_facout), .Cin(s5_522_facout), .S(s6_530_fas), .Cout(s6_530_facout));
full_adder s6_53fa1 ( .A(s5_530_fas), .B(s5_531_fas), .Cin(s5_532_fas), .S(s6_531_fas), .Cout(s6_531_facout));
full_adder s6_54fa0 ( .A(s5_530_facout), .B(s5_531_facout), .Cin(s5_532_facout), .S(s6_540_fas), .Cout(s6_540_facout));
full_adder s6_54fa1 ( .A(s5_540_fas), .B(s5_541_fas), .Cin(s5_542_fas), .S(s6_541_fas), .Cout(s6_541_facout));
full_adder s6_55fa0 ( .A(s5_540_facout), .B(s5_541_facout), .Cin(s5_542_facout), .S(s6_550_fas), .Cout(s6_550_facout));
full_adder s6_55fa1 ( .A(s5_550_fas), .B(s5_551_fas), .Cin(s5_552_fas), .S(s6_551_fas), .Cout(s6_551_facout));
full_adder s6_56fa0 ( .A(ps_5625), .B(s5_550_facout), .Cin(s5_551_facout), .S(s6_560_fas), .Cout(s6_560_facout));
full_adder s6_56fa1 ( .A(s5_552_facout), .B(s5_560_fas), .Cin(s5_561_fas), .S(s6_561_fas), .Cout(s6_561_facout));
full_adder s6_57fa0 ( .A(ps_5728), .B(ps_5727), .Cin(ps_5726), .S(s6_570_fas), .Cout(s6_570_facout));
full_adder s6_57fa1 ( .A(s5_560_facout), .B(s5_561_facout), .Cin(s5_570_fas), .S(s6_571_fas), .Cout(s6_571_facout));
full_adder s6_58fa0 ( .A(ps_5831), .B(ps_5830), .Cin(ps_5829), .S(s6_580_fas), .Cout(s6_580_facout));
full_adder s6_58fa1 ( .A(ps_5828), .B(ps_5827), .Cin(s5_570_facout), .S(s6_581_fas), .Cout(s6_581_facout));
full_adder s6_59fa0 ( .A(ps_5931), .B(ps_5930), .Cin(ps_5929), .S(s6_590_fas), .Cout(s6_590_facout));
logic s7_30_hacout, s7_30_has, s7_40_facout, s7_40_fas, s7_50_facout, s7_50_fas, s7_60_facout, s7_60_fas, s7_70_facout, s7_70_fas, s7_80_facout, s7_80_fas, s7_90_facout, s7_90_fas, s7_100_facout, s7_100_fas, s7_110_facout, s7_110_fas, s7_120_facout, s7_120_fas, s7_130_facout, s7_130_fas, s7_140_facout, s7_140_fas, s7_150_facout, s7_150_fas, s7_160_facout, s7_160_fas, s7_170_facout, s7_170_fas, s7_180_facout, s7_180_fas, s7_190_facout, s7_190_fas, s7_200_facout, s7_200_fas, s7_210_facout, s7_210_fas, s7_220_facout, s7_220_fas, s7_230_facout, s7_230_fas, s7_240_facout, s7_240_fas, s7_250_facout, s7_250_fas, s7_260_facout, s7_260_fas, s7_270_facout, s7_270_fas, s7_280_facout, s7_280_fas, s7_290_facout, s7_290_fas, s7_300_facout, s7_300_fas, s7_310_facout, s7_310_fas, s7_320_facout, s7_320_fas, s7_330_facout, s7_330_fas, s7_340_facout, s7_340_fas, s7_350_facout, s7_350_fas, s7_360_facout, s7_360_fas, s7_370_facout, s7_370_fas, s7_380_facout, s7_380_fas, s7_390_facout, s7_390_fas, s7_400_facout, s7_400_fas, s7_410_facout, s7_410_fas, s7_420_facout, s7_420_fas, s7_430_facout, s7_430_fas, s7_440_facout, s7_440_fas, s7_450_facout, s7_450_fas, s7_460_facout, s7_460_fas, s7_470_facout, s7_470_fas, s7_480_facout, s7_480_fas, s7_490_facout, s7_490_fas, s7_500_facout, s7_500_fas, s7_510_facout, s7_510_fas, s7_520_facout, s7_520_fas, s7_530_facout, s7_530_fas, s7_540_facout, s7_540_fas, s7_550_facout, s7_550_fas, s7_560_facout, s7_560_fas, s7_570_facout, s7_570_fas, s7_580_facout, s7_580_fas, s7_590_facout, s7_590_fas, s7_600_facout, s7_600_fas;
/* ========================= Stage 7 ========================= */
half_adder s7_3ha0 ( .A(ps_33), .B(ps_32), .S(s7_30_has), .Cout(s7_30_hacout));
full_adder s7_4fa0 ( .A(ps_42), .B(ps_41), .Cin(ps_40), .S(s7_40_fas), .Cout(s7_40_facout));
full_adder s7_5fa0 ( .A(ps_50), .B(s6_40_hacout), .Cin(s6_50_fas), .S(s7_50_fas), .Cout(s7_50_facout));
full_adder s7_6fa0 ( .A(s6_50_facout), .B(s6_50_hacout), .Cin(s6_60_fas), .S(s7_60_fas), .Cout(s7_60_facout));
full_adder s7_7fa0 ( .A(s6_60_facout), .B(s6_61_facout), .Cin(s6_70_fas), .S(s7_70_fas), .Cout(s7_70_facout));
full_adder s7_8fa0 ( .A(s6_70_facout), .B(s6_71_facout), .Cin(s6_80_fas), .S(s7_80_fas), .Cout(s7_80_facout));
full_adder s7_9fa0 ( .A(s6_80_facout), .B(s6_81_facout), .Cin(s6_90_fas), .S(s7_90_fas), .Cout(s7_90_facout));
full_adder s7_10fa0 ( .A(s6_90_facout), .B(s6_91_facout), .Cin(s6_100_fas), .S(s7_100_fas), .Cout(s7_100_facout));
full_adder s7_11fa0 ( .A(s6_100_facout), .B(s6_101_facout), .Cin(s6_110_fas), .S(s7_110_fas), .Cout(s7_110_facout));
full_adder s7_12fa0 ( .A(s6_110_facout), .B(s6_111_facout), .Cin(s6_120_fas), .S(s7_120_fas), .Cout(s7_120_facout));
full_adder s7_13fa0 ( .A(s6_120_facout), .B(s6_121_facout), .Cin(s6_130_fas), .S(s7_130_fas), .Cout(s7_130_facout));
full_adder s7_14fa0 ( .A(s6_130_facout), .B(s6_131_facout), .Cin(s6_140_fas), .S(s7_140_fas), .Cout(s7_140_facout));
full_adder s7_15fa0 ( .A(s6_140_facout), .B(s6_141_facout), .Cin(s6_150_fas), .S(s7_150_fas), .Cout(s7_150_facout));
full_adder s7_16fa0 ( .A(s6_150_facout), .B(s6_151_facout), .Cin(s6_160_fas), .S(s7_160_fas), .Cout(s7_160_facout));
full_adder s7_17fa0 ( .A(s6_160_facout), .B(s6_161_facout), .Cin(s6_170_fas), .S(s7_170_fas), .Cout(s7_170_facout));
full_adder s7_18fa0 ( .A(s6_170_facout), .B(s6_171_facout), .Cin(s6_180_fas), .S(s7_180_fas), .Cout(s7_180_facout));
full_adder s7_19fa0 ( .A(s6_180_facout), .B(s6_181_facout), .Cin(s6_190_fas), .S(s7_190_fas), .Cout(s7_190_facout));
full_adder s7_20fa0 ( .A(s6_190_facout), .B(s6_191_facout), .Cin(s6_200_fas), .S(s7_200_fas), .Cout(s7_200_facout));
full_adder s7_21fa0 ( .A(s6_200_facout), .B(s6_201_facout), .Cin(s6_210_fas), .S(s7_210_fas), .Cout(s7_210_facout));
full_adder s7_22fa0 ( .A(s6_210_facout), .B(s6_211_facout), .Cin(s6_220_fas), .S(s7_220_fas), .Cout(s7_220_facout));
full_adder s7_23fa0 ( .A(s6_220_facout), .B(s6_221_facout), .Cin(s6_230_fas), .S(s7_230_fas), .Cout(s7_230_facout));
full_adder s7_24fa0 ( .A(s6_230_facout), .B(s6_231_facout), .Cin(s6_240_fas), .S(s7_240_fas), .Cout(s7_240_facout));
full_adder s7_25fa0 ( .A(s6_240_facout), .B(s6_241_facout), .Cin(s6_250_fas), .S(s7_250_fas), .Cout(s7_250_facout));
full_adder s7_26fa0 ( .A(s6_250_facout), .B(s6_251_facout), .Cin(s6_260_fas), .S(s7_260_fas), .Cout(s7_260_facout));
full_adder s7_27fa0 ( .A(s6_260_facout), .B(s6_261_facout), .Cin(s6_270_fas), .S(s7_270_fas), .Cout(s7_270_facout));
full_adder s7_28fa0 ( .A(s6_270_facout), .B(s6_271_facout), .Cin(s6_280_fas), .S(s7_280_fas), .Cout(s7_280_facout));
full_adder s7_29fa0 ( .A(s6_280_facout), .B(s6_281_facout), .Cin(s6_290_fas), .S(s7_290_fas), .Cout(s7_290_facout));
full_adder s7_30fa0 ( .A(s6_290_facout), .B(s6_291_facout), .Cin(s6_300_fas), .S(s7_300_fas), .Cout(s7_300_facout));
full_adder s7_31fa0 ( .A(s6_300_facout), .B(s6_301_facout), .Cin(s6_310_fas), .S(s7_310_fas), .Cout(s7_310_facout));
full_adder s7_32fa0 ( .A(s6_310_facout), .B(s6_311_facout), .Cin(s6_320_fas), .S(s7_320_fas), .Cout(s7_320_facout));
full_adder s7_33fa0 ( .A(s6_320_facout), .B(s6_321_facout), .Cin(s6_330_fas), .S(s7_330_fas), .Cout(s7_330_facout));
full_adder s7_34fa0 ( .A(s6_330_facout), .B(s6_331_facout), .Cin(s6_340_fas), .S(s7_340_fas), .Cout(s7_340_facout));
full_adder s7_35fa0 ( .A(s6_340_facout), .B(s6_341_facout), .Cin(s6_350_fas), .S(s7_350_fas), .Cout(s7_350_facout));
full_adder s7_36fa0 ( .A(s6_350_facout), .B(s6_351_facout), .Cin(s6_360_fas), .S(s7_360_fas), .Cout(s7_360_facout));
full_adder s7_37fa0 ( .A(s6_360_facout), .B(s6_361_facout), .Cin(s6_370_fas), .S(s7_370_fas), .Cout(s7_370_facout));
full_adder s7_38fa0 ( .A(s6_370_facout), .B(s6_371_facout), .Cin(s6_380_fas), .S(s7_380_fas), .Cout(s7_380_facout));
full_adder s7_39fa0 ( .A(s6_380_facout), .B(s6_381_facout), .Cin(s6_390_fas), .S(s7_390_fas), .Cout(s7_390_facout));
full_adder s7_40fa0 ( .A(s6_390_facout), .B(s6_391_facout), .Cin(s6_400_fas), .S(s7_400_fas), .Cout(s7_400_facout));
full_adder s7_41fa0 ( .A(s6_400_facout), .B(s6_401_facout), .Cin(s6_410_fas), .S(s7_410_fas), .Cout(s7_410_facout));
full_adder s7_42fa0 ( .A(s6_410_facout), .B(s6_411_facout), .Cin(s6_420_fas), .S(s7_420_fas), .Cout(s7_420_facout));
full_adder s7_43fa0 ( .A(s6_420_facout), .B(s6_421_facout), .Cin(s6_430_fas), .S(s7_430_fas), .Cout(s7_430_facout));
full_adder s7_44fa0 ( .A(s6_430_facout), .B(s6_431_facout), .Cin(s6_440_fas), .S(s7_440_fas), .Cout(s7_440_facout));
full_adder s7_45fa0 ( .A(s6_440_facout), .B(s6_441_facout), .Cin(s6_450_fas), .S(s7_450_fas), .Cout(s7_450_facout));
full_adder s7_46fa0 ( .A(s6_450_facout), .B(s6_451_facout), .Cin(s6_460_fas), .S(s7_460_fas), .Cout(s7_460_facout));
full_adder s7_47fa0 ( .A(s6_460_facout), .B(s6_461_facout), .Cin(s6_470_fas), .S(s7_470_fas), .Cout(s7_470_facout));
full_adder s7_48fa0 ( .A(s6_470_facout), .B(s6_471_facout), .Cin(s6_480_fas), .S(s7_480_fas), .Cout(s7_480_facout));
full_adder s7_49fa0 ( .A(s6_480_facout), .B(s6_481_facout), .Cin(s6_490_fas), .S(s7_490_fas), .Cout(s7_490_facout));
full_adder s7_50fa0 ( .A(s6_490_facout), .B(s6_491_facout), .Cin(s6_500_fas), .S(s7_500_fas), .Cout(s7_500_facout));
full_adder s7_51fa0 ( .A(s6_500_facout), .B(s6_501_facout), .Cin(s6_510_fas), .S(s7_510_fas), .Cout(s7_510_facout));
full_adder s7_52fa0 ( .A(s6_510_facout), .B(s6_511_facout), .Cin(s6_520_fas), .S(s7_520_fas), .Cout(s7_520_facout));
full_adder s7_53fa0 ( .A(s6_520_facout), .B(s6_521_facout), .Cin(s6_530_fas), .S(s7_530_fas), .Cout(s7_530_facout));
full_adder s7_54fa0 ( .A(s6_530_facout), .B(s6_531_facout), .Cin(s6_540_fas), .S(s7_540_fas), .Cout(s7_540_facout));
full_adder s7_55fa0 ( .A(s6_540_facout), .B(s6_541_facout), .Cin(s6_550_fas), .S(s7_550_fas), .Cout(s7_550_facout));
full_adder s7_56fa0 ( .A(s6_550_facout), .B(s6_551_facout), .Cin(s6_560_fas), .S(s7_560_fas), .Cout(s7_560_facout));
full_adder s7_57fa0 ( .A(s6_560_facout), .B(s6_561_facout), .Cin(s6_570_fas), .S(s7_570_fas), .Cout(s7_570_facout));
full_adder s7_58fa0 ( .A(s6_570_facout), .B(s6_571_facout), .Cin(s6_580_fas), .S(s7_580_fas), .Cout(s7_580_facout));
full_adder s7_59fa0 ( .A(ps_5928), .B(s6_580_facout), .Cin(s6_581_facout), .S(s7_590_fas), .Cout(s7_590_facout));
full_adder s7_60fa0 ( .A(ps_6031), .B(ps_6030), .Cin(ps_6029), .S(s7_600_fas), .Cout(s7_600_facout));
logic s8_20_hacout, s8_20_has, s8_30_facout, s8_30_fas, s8_40_facout, s8_40_fas, s8_50_facout, s8_50_fas, s8_60_facout, s8_60_fas, s8_70_facout, s8_70_fas, s8_80_facout, s8_80_fas, s8_90_facout, s8_90_fas, s8_100_facout, s8_100_fas, s8_110_facout, s8_110_fas, s8_120_facout, s8_120_fas, s8_130_facout, s8_130_fas, s8_140_facout, s8_140_fas, s8_150_facout, s8_150_fas, s8_160_facout, s8_160_fas, s8_170_facout, s8_170_fas, s8_180_facout, s8_180_fas, s8_190_facout, s8_190_fas, s8_200_facout, s8_200_fas, s8_210_facout, s8_210_fas, s8_220_facout, s8_220_fas, s8_230_facout, s8_230_fas, s8_240_facout, s8_240_fas, s8_250_facout, s8_250_fas, s8_260_facout, s8_260_fas, s8_270_facout, s8_270_fas, s8_280_facout, s8_280_fas, s8_290_facout, s8_290_fas, s8_300_facout, s8_300_fas, s8_310_facout, s8_310_fas, s8_320_facout, s8_320_fas, s8_330_facout, s8_330_fas, s8_340_facout, s8_340_fas, s8_350_facout, s8_350_fas, s8_360_facout, s8_360_fas, s8_370_facout, s8_370_fas, s8_380_facout, s8_380_fas, s8_390_facout, s8_390_fas, s8_400_facout, s8_400_fas, s8_410_facout, s8_410_fas, s8_420_facout, s8_420_fas, s8_430_facout, s8_430_fas, s8_440_facout, s8_440_fas, s8_450_facout, s8_450_fas, s8_460_facout, s8_460_fas, s8_470_facout, s8_470_fas, s8_480_facout, s8_480_fas, s8_490_facout, s8_490_fas, s8_500_facout, s8_500_fas, s8_510_facout, s8_510_fas, s8_520_facout, s8_520_fas, s8_530_facout, s8_530_fas, s8_540_facout, s8_540_fas, s8_550_facout, s8_550_fas, s8_560_facout, s8_560_fas, s8_570_facout, s8_570_fas, s8_580_facout, s8_580_fas, s8_590_facout, s8_590_fas, s8_600_facout, s8_600_fas, s8_610_facout, s8_610_fas;
/* ========================= Stage 8 ========================= */
half_adder s8_2ha0 ( .A(ps_22), .B(ps_21), .S(s8_20_has), .Cout(s8_20_hacout));
full_adder s8_3fa0 ( .A(ps_31), .B(ps_30), .Cin(s7_30_has), .S(s8_30_fas), .Cout(s8_30_facout));
full_adder s8_4fa0 ( .A(s6_40_has), .B(s7_30_hacout), .Cin(s7_40_fas), .S(s8_40_fas), .Cout(s8_40_facout));
full_adder s8_5fa0 ( .A(s6_50_has), .B(s7_40_facout), .Cin(s7_50_fas), .S(s8_50_fas), .Cout(s8_50_facout));
full_adder s8_6fa0 ( .A(s6_61_fas), .B(s7_50_facout), .Cin(s7_60_fas), .S(s8_60_fas), .Cout(s8_60_facout));
full_adder s8_7fa0 ( .A(s6_71_fas), .B(s7_60_facout), .Cin(s7_70_fas), .S(s8_70_fas), .Cout(s8_70_facout));
full_adder s8_8fa0 ( .A(s6_81_fas), .B(s7_70_facout), .Cin(s7_80_fas), .S(s8_80_fas), .Cout(s8_80_facout));
full_adder s8_9fa0 ( .A(s6_91_fas), .B(s7_80_facout), .Cin(s7_90_fas), .S(s8_90_fas), .Cout(s8_90_facout));
full_adder s8_10fa0 ( .A(s6_101_fas), .B(s7_90_facout), .Cin(s7_100_fas), .S(s8_100_fas), .Cout(s8_100_facout));
full_adder s8_11fa0 ( .A(s6_111_fas), .B(s7_100_facout), .Cin(s7_110_fas), .S(s8_110_fas), .Cout(s8_110_facout));
full_adder s8_12fa0 ( .A(s6_121_fas), .B(s7_110_facout), .Cin(s7_120_fas), .S(s8_120_fas), .Cout(s8_120_facout));
full_adder s8_13fa0 ( .A(s6_131_fas), .B(s7_120_facout), .Cin(s7_130_fas), .S(s8_130_fas), .Cout(s8_130_facout));
full_adder s8_14fa0 ( .A(s6_141_fas), .B(s7_130_facout), .Cin(s7_140_fas), .S(s8_140_fas), .Cout(s8_140_facout));
full_adder s8_15fa0 ( .A(s6_151_fas), .B(s7_140_facout), .Cin(s7_150_fas), .S(s8_150_fas), .Cout(s8_150_facout));
full_adder s8_16fa0 ( .A(s6_161_fas), .B(s7_150_facout), .Cin(s7_160_fas), .S(s8_160_fas), .Cout(s8_160_facout));
full_adder s8_17fa0 ( .A(s6_171_fas), .B(s7_160_facout), .Cin(s7_170_fas), .S(s8_170_fas), .Cout(s8_170_facout));
full_adder s8_18fa0 ( .A(s6_181_fas), .B(s7_170_facout), .Cin(s7_180_fas), .S(s8_180_fas), .Cout(s8_180_facout));
full_adder s8_19fa0 ( .A(s6_191_fas), .B(s7_180_facout), .Cin(s7_190_fas), .S(s8_190_fas), .Cout(s8_190_facout));
full_adder s8_20fa0 ( .A(s6_201_fas), .B(s7_190_facout), .Cin(s7_200_fas), .S(s8_200_fas), .Cout(s8_200_facout));
full_adder s8_21fa0 ( .A(s6_211_fas), .B(s7_200_facout), .Cin(s7_210_fas), .S(s8_210_fas), .Cout(s8_210_facout));
full_adder s8_22fa0 ( .A(s6_221_fas), .B(s7_210_facout), .Cin(s7_220_fas), .S(s8_220_fas), .Cout(s8_220_facout));
full_adder s8_23fa0 ( .A(s6_231_fas), .B(s7_220_facout), .Cin(s7_230_fas), .S(s8_230_fas), .Cout(s8_230_facout));
full_adder s8_24fa0 ( .A(s6_241_fas), .B(s7_230_facout), .Cin(s7_240_fas), .S(s8_240_fas), .Cout(s8_240_facout));
full_adder s8_25fa0 ( .A(s6_251_fas), .B(s7_240_facout), .Cin(s7_250_fas), .S(s8_250_fas), .Cout(s8_250_facout));
full_adder s8_26fa0 ( .A(s6_261_fas), .B(s7_250_facout), .Cin(s7_260_fas), .S(s8_260_fas), .Cout(s8_260_facout));
full_adder s8_27fa0 ( .A(s6_271_fas), .B(s7_260_facout), .Cin(s7_270_fas), .S(s8_270_fas), .Cout(s8_270_facout));
full_adder s8_28fa0 ( .A(s6_281_fas), .B(s7_270_facout), .Cin(s7_280_fas), .S(s8_280_fas), .Cout(s8_280_facout));
full_adder s8_29fa0 ( .A(s6_291_fas), .B(s7_280_facout), .Cin(s7_290_fas), .S(s8_290_fas), .Cout(s8_290_facout));
full_adder s8_30fa0 ( .A(s6_301_fas), .B(s7_290_facout), .Cin(s7_300_fas), .S(s8_300_fas), .Cout(s8_300_facout));
full_adder s8_31fa0 ( .A(s6_311_fas), .B(s7_300_facout), .Cin(s7_310_fas), .S(s8_310_fas), .Cout(s8_310_facout));
full_adder s8_32fa0 ( .A(s6_321_fas), .B(s7_310_facout), .Cin(s7_320_fas), .S(s8_320_fas), .Cout(s8_320_facout));
full_adder s8_33fa0 ( .A(s6_331_fas), .B(s7_320_facout), .Cin(s7_330_fas), .S(s8_330_fas), .Cout(s8_330_facout));
full_adder s8_34fa0 ( .A(s6_341_fas), .B(s7_330_facout), .Cin(s7_340_fas), .S(s8_340_fas), .Cout(s8_340_facout));
full_adder s8_35fa0 ( .A(s6_351_fas), .B(s7_340_facout), .Cin(s7_350_fas), .S(s8_350_fas), .Cout(s8_350_facout));
full_adder s8_36fa0 ( .A(s6_361_fas), .B(s7_350_facout), .Cin(s7_360_fas), .S(s8_360_fas), .Cout(s8_360_facout));
full_adder s8_37fa0 ( .A(s6_371_fas), .B(s7_360_facout), .Cin(s7_370_fas), .S(s8_370_fas), .Cout(s8_370_facout));
full_adder s8_38fa0 ( .A(s6_381_fas), .B(s7_370_facout), .Cin(s7_380_fas), .S(s8_380_fas), .Cout(s8_380_facout));
full_adder s8_39fa0 ( .A(s6_391_fas), .B(s7_380_facout), .Cin(s7_390_fas), .S(s8_390_fas), .Cout(s8_390_facout));
full_adder s8_40fa0 ( .A(s6_401_fas), .B(s7_390_facout), .Cin(s7_400_fas), .S(s8_400_fas), .Cout(s8_400_facout));
full_adder s8_41fa0 ( .A(s6_411_fas), .B(s7_400_facout), .Cin(s7_410_fas), .S(s8_410_fas), .Cout(s8_410_facout));
full_adder s8_42fa0 ( .A(s6_421_fas), .B(s7_410_facout), .Cin(s7_420_fas), .S(s8_420_fas), .Cout(s8_420_facout));
full_adder s8_43fa0 ( .A(s6_431_fas), .B(s7_420_facout), .Cin(s7_430_fas), .S(s8_430_fas), .Cout(s8_430_facout));
full_adder s8_44fa0 ( .A(s6_441_fas), .B(s7_430_facout), .Cin(s7_440_fas), .S(s8_440_fas), .Cout(s8_440_facout));
full_adder s8_45fa0 ( .A(s6_451_fas), .B(s7_440_facout), .Cin(s7_450_fas), .S(s8_450_fas), .Cout(s8_450_facout));
full_adder s8_46fa0 ( .A(s6_461_fas), .B(s7_450_facout), .Cin(s7_460_fas), .S(s8_460_fas), .Cout(s8_460_facout));
full_adder s8_47fa0 ( .A(s6_471_fas), .B(s7_460_facout), .Cin(s7_470_fas), .S(s8_470_fas), .Cout(s8_470_facout));
full_adder s8_48fa0 ( .A(s6_481_fas), .B(s7_470_facout), .Cin(s7_480_fas), .S(s8_480_fas), .Cout(s8_480_facout));
full_adder s8_49fa0 ( .A(s6_491_fas), .B(s7_480_facout), .Cin(s7_490_fas), .S(s8_490_fas), .Cout(s8_490_facout));
full_adder s8_50fa0 ( .A(s6_501_fas), .B(s7_490_facout), .Cin(s7_500_fas), .S(s8_500_fas), .Cout(s8_500_facout));
full_adder s8_51fa0 ( .A(s6_511_fas), .B(s7_500_facout), .Cin(s7_510_fas), .S(s8_510_fas), .Cout(s8_510_facout));
full_adder s8_52fa0 ( .A(s6_521_fas), .B(s7_510_facout), .Cin(s7_520_fas), .S(s8_520_fas), .Cout(s8_520_facout));
full_adder s8_53fa0 ( .A(s6_531_fas), .B(s7_520_facout), .Cin(s7_530_fas), .S(s8_530_fas), .Cout(s8_530_facout));
full_adder s8_54fa0 ( .A(s6_541_fas), .B(s7_530_facout), .Cin(s7_540_fas), .S(s8_540_fas), .Cout(s8_540_facout));
full_adder s8_55fa0 ( .A(s6_551_fas), .B(s7_540_facout), .Cin(s7_550_fas), .S(s8_550_fas), .Cout(s8_550_facout));
full_adder s8_56fa0 ( .A(s6_561_fas), .B(s7_550_facout), .Cin(s7_560_fas), .S(s8_560_fas), .Cout(s8_560_facout));
full_adder s8_57fa0 ( .A(s6_571_fas), .B(s7_560_facout), .Cin(s7_570_fas), .S(s8_570_fas), .Cout(s8_570_facout));
full_adder s8_58fa0 ( .A(s6_581_fas), .B(s7_570_facout), .Cin(s7_580_fas), .S(s8_580_fas), .Cout(s8_580_facout));
full_adder s8_59fa0 ( .A(s6_590_fas), .B(s7_580_facout), .Cin(s7_590_fas), .S(s8_590_fas), .Cout(s8_590_facout));
full_adder s8_60fa0 ( .A(s6_590_facout), .B(s7_590_facout), .Cin(s7_600_fas), .S(s8_600_fas), .Cout(s8_600_facout));
full_adder s8_61fa0 ( .A(ps_6131), .B(ps_6130), .Cin(s7_600_facout), .S(s8_610_fas), .Cout(s8_610_facout));
logic [63:0] op1, op2;
assign op1[0] = ps_00;
assign op2[0] = '0;
assign op1[1] = ps_11;
assign op2[1] = ps_10;
assign op1[2] = ps_20;
assign op2[2] = s8_20_has;
assign op1[3] = s8_20_hacout;
assign op2[3] = s8_30_fas;
assign op1[4] = s8_30_facout;
assign op2[4] = s8_40_fas;
assign op1[5] = s8_40_facout;
assign op2[5] = s8_50_fas;
assign op1[6] = s8_50_facout;
assign op2[6] = s8_60_fas;
assign op1[7] = s8_60_facout;
assign op2[7] = s8_70_fas;
assign op1[8] = s8_70_facout;
assign op2[8] = s8_80_fas;
assign op1[9] = s8_80_facout;
assign op2[9] = s8_90_fas;
assign op1[10] = s8_90_facout;
assign op2[10] = s8_100_fas;
assign op1[11] = s8_100_facout;
assign op2[11] = s8_110_fas;
assign op1[12] = s8_110_facout;
assign op2[12] = s8_120_fas;
assign op1[13] = s8_120_facout;
assign op2[13] = s8_130_fas;
assign op1[14] = s8_130_facout;
assign op2[14] = s8_140_fas;
assign op1[15] = s8_140_facout;
assign op2[15] = s8_150_fas;
assign op1[16] = s8_150_facout;
assign op2[16] = s8_160_fas;
assign op1[17] = s8_160_facout;
assign op2[17] = s8_170_fas;
assign op1[18] = s8_170_facout;
assign op2[18] = s8_180_fas;
assign op1[19] = s8_180_facout;
assign op2[19] = s8_190_fas;
assign op1[20] = s8_190_facout;
assign op2[20] = s8_200_fas;
assign op1[21] = s8_200_facout;
assign op2[21] = s8_210_fas;
assign op1[22] = s8_210_facout;
assign op2[22] = s8_220_fas;
assign op1[23] = s8_220_facout;
assign op2[23] = s8_230_fas;
assign op1[24] = s8_230_facout;
assign op2[24] = s8_240_fas;
assign op1[25] = s8_240_facout;
assign op2[25] = s8_250_fas;
assign op1[26] = s8_250_facout;
assign op2[26] = s8_260_fas;
assign op1[27] = s8_260_facout;
assign op2[27] = s8_270_fas;
assign op1[28] = s8_270_facout;
assign op2[28] = s8_280_fas;
assign op1[29] = s8_280_facout;
assign op2[29] = s8_290_fas;
assign op1[30] = s8_290_facout;
assign op2[30] = s8_300_fas;
assign op1[31] = s8_300_facout;
assign op2[31] = s8_310_fas;
assign op1[32] = s8_310_facout;
assign op2[32] = s8_320_fas;
assign op1[33] = s8_320_facout;
assign op2[33] = s8_330_fas;
assign op1[34] = s8_330_facout;
assign op2[34] = s8_340_fas;
assign op1[35] = s8_340_facout;
assign op2[35] = s8_350_fas;
assign op1[36] = s8_350_facout;
assign op2[36] = s8_360_fas;
assign op1[37] = s8_360_facout;
assign op2[37] = s8_370_fas;
assign op1[38] = s8_370_facout;
assign op2[38] = s8_380_fas;
assign op1[39] = s8_380_facout;
assign op2[39] = s8_390_fas;
assign op1[40] = s8_390_facout;
assign op2[40] = s8_400_fas;
assign op1[41] = s8_400_facout;
assign op2[41] = s8_410_fas;
assign op1[42] = s8_410_facout;
assign op2[42] = s8_420_fas;
assign op1[43] = s8_420_facout;
assign op2[43] = s8_430_fas;
assign op1[44] = s8_430_facout;
assign op2[44] = s8_440_fas;
assign op1[45] = s8_440_facout;
assign op2[45] = s8_450_fas;
assign op1[46] = s8_450_facout;
assign op2[46] = s8_460_fas;
assign op1[47] = s8_460_facout;
assign op2[47] = s8_470_fas;
assign op1[48] = s8_470_facout;
assign op2[48] = s8_480_fas;
assign op1[49] = s8_480_facout;
assign op2[49] = s8_490_fas;
assign op1[50] = s8_490_facout;
assign op2[50] = s8_500_fas;
assign op1[51] = s8_500_facout;
assign op2[51] = s8_510_fas;
assign op1[52] = s8_510_facout;
assign op2[52] = s8_520_fas;
assign op1[53] = s8_520_facout;
assign op2[53] = s8_530_fas;
assign op1[54] = s8_530_facout;
assign op2[54] = s8_540_fas;
assign op1[55] = s8_540_facout;
assign op2[55] = s8_550_fas;
assign op1[56] = s8_550_facout;
assign op2[56] = s8_560_fas;
assign op1[57] = s8_560_facout;
assign op2[57] = s8_570_fas;
assign op1[58] = s8_570_facout;
assign op2[58] = s8_580_fas;
assign op1[59] = s8_580_facout;
assign op2[59] = s8_590_fas;
assign op1[60] = s8_590_facout;
assign op2[60] = s8_600_fas;
assign op1[61] = s8_600_facout;
assign op2[61] = s8_610_fas;
assign op1[62] = ps_6231;
assign op2[62] = s8_610_facout;
assign op1[63] = '0;
assign op2[63] = '0;
assign pre_result_in = op1 + op2;

endmodule